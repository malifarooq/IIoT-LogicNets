module layer1 (input [1023:0] M0, output [171:0] M1);

wire [11:0] layer1_N0_wire = {M0[999], M0[998], M0[965], M0[964], M0[523], M0[522], M0[451], M0[450], M0[195], M0[194], M0[97], M0[96]};
layer1_N0 layer1_N0_inst (.M0(layer1_N0_wire), .M1(M1[1:0]));

wire [11:0] layer1_N1_wire = {M0[963], M0[962], M0[621], M0[620], M0[615], M0[614], M0[481], M0[480], M0[367], M0[366], M0[55], M0[54]};
layer1_N1 layer1_N1_inst (.M0(layer1_N1_wire), .M1(M1[3:2]));

wire [11:0] layer1_N2_wire = {M0[999], M0[998], M0[985], M0[984], M0[665], M0[664], M0[507], M0[506], M0[323], M0[322], M0[189], M0[188]};
layer1_N2 layer1_N2_inst (.M0(layer1_N2_wire), .M1(M1[5:4]));

wire [11:0] layer1_N3_wire = {M0[937], M0[936], M0[931], M0[930], M0[671], M0[670], M0[509], M0[508], M0[369], M0[368], M0[253], M0[252]};
layer1_N3 layer1_N3_inst (.M0(layer1_N3_wire), .M1(M1[7:6]));

wire [11:0] layer1_N4_wire = {M0[901], M0[900], M0[549], M0[548], M0[399], M0[398], M0[367], M0[366], M0[99], M0[98], M0[13], M0[12]};
layer1_N4 layer1_N4_inst (.M0(layer1_N4_wire), .M1(M1[9:8]));

wire [11:0] layer1_N5_wire = {M0[991], M0[990], M0[825], M0[824], M0[695], M0[694], M0[689], M0[688], M0[247], M0[246], M0[99], M0[98]};
layer1_N5 layer1_N5_inst (.M0(layer1_N5_wire), .M1(M1[11:10]));

wire [11:0] layer1_N6_wire = {M0[825], M0[824], M0[685], M0[684], M0[491], M0[490], M0[195], M0[194], M0[165], M0[164], M0[29], M0[28]};
layer1_N6 layer1_N6_inst (.M0(layer1_N6_wire), .M1(M1[13:12]));

wire [11:0] layer1_N7_wire = {M0[961], M0[960], M0[867], M0[866], M0[809], M0[808], M0[287], M0[286], M0[283], M0[282], M0[3], M0[2]};
layer1_N7 layer1_N7_inst (.M0(layer1_N7_wire), .M1(M1[15:14]));

wire [11:0] layer1_N8_wire = {M0[1001], M0[1000], M0[605], M0[604], M0[335], M0[334], M0[307], M0[306], M0[255], M0[254], M0[193], M0[192]};
layer1_N8 layer1_N8_inst (.M0(layer1_N8_wire), .M1(M1[17:16]));

wire [11:0] layer1_N9_wire = {M0[819], M0[818], M0[811], M0[810], M0[739], M0[738], M0[489], M0[488], M0[405], M0[404], M0[113], M0[112]};
layer1_N9 layer1_N9_inst (.M0(layer1_N9_wire), .M1(M1[19:18]));

wire [11:0] layer1_N10_wire = {M0[929], M0[928], M0[757], M0[756], M0[635], M0[634], M0[297], M0[296], M0[227], M0[226], M0[61], M0[60]};
layer1_N10 layer1_N10_inst (.M0(layer1_N10_wire), .M1(M1[21:20]));

wire [11:0] layer1_N11_wire = {M0[677], M0[676], M0[675], M0[674], M0[519], M0[518], M0[327], M0[326], M0[289], M0[288], M0[215], M0[214]};
layer1_N11 layer1_N11_inst (.M0(layer1_N11_wire), .M1(M1[23:22]));

wire [11:0] layer1_N12_wire = {M0[957], M0[956], M0[927], M0[926], M0[421], M0[420], M0[387], M0[386], M0[269], M0[268], M0[139], M0[138]};
layer1_N12 layer1_N12_inst (.M0(layer1_N12_wire), .M1(M1[25:24]));

wire [11:0] layer1_N13_wire = {M0[771], M0[770], M0[599], M0[598], M0[433], M0[432], M0[429], M0[428], M0[257], M0[256], M0[47], M0[46]};
layer1_N13 layer1_N13_inst (.M0(layer1_N13_wire), .M1(M1[27:26]));

wire [11:0] layer1_N14_wire = {M0[787], M0[786], M0[723], M0[722], M0[675], M0[674], M0[409], M0[408], M0[165], M0[164], M0[55], M0[54]};
layer1_N14 layer1_N14_inst (.M0(layer1_N14_wire), .M1(M1[29:28]));

wire [11:0] layer1_N15_wire = {M0[1023], M0[1022], M0[869], M0[868], M0[695], M0[694], M0[415], M0[414], M0[241], M0[240], M0[167], M0[166]};
layer1_N15 layer1_N15_inst (.M0(layer1_N15_wire), .M1(M1[31:30]));

wire [11:0] layer1_N16_wire = {M0[799], M0[798], M0[603], M0[602], M0[529], M0[528], M0[475], M0[474], M0[297], M0[296], M0[115], M0[114]};
layer1_N16 layer1_N16_inst (.M0(layer1_N16_wire), .M1(M1[33:32]));

wire [11:0] layer1_N17_wire = {M0[1003], M0[1002], M0[953], M0[952], M0[925], M0[924], M0[679], M0[678], M0[403], M0[402], M0[103], M0[102]};
layer1_N17 layer1_N17_inst (.M0(layer1_N17_wire), .M1(M1[35:34]));

wire [11:0] layer1_N18_wire = {M0[843], M0[842], M0[835], M0[834], M0[787], M0[786], M0[521], M0[520], M0[441], M0[440], M0[335], M0[334]};
layer1_N18 layer1_N18_inst (.M0(layer1_N18_wire), .M1(M1[37:36]));

wire [11:0] layer1_N19_wire = {M0[1005], M0[1004], M0[931], M0[930], M0[737], M0[736], M0[593], M0[592], M0[385], M0[384], M0[199], M0[198]};
layer1_N19 layer1_N19_inst (.M0(layer1_N19_wire), .M1(M1[39:38]));

wire [11:0] layer1_N20_wire = {M0[837], M0[836], M0[679], M0[678], M0[673], M0[672], M0[345], M0[344], M0[207], M0[206], M0[205], M0[204]};
layer1_N20 layer1_N20_inst (.M0(layer1_N20_wire), .M1(M1[41:40]));

wire [11:0] layer1_N21_wire = {M0[957], M0[956], M0[921], M0[920], M0[665], M0[664], M0[609], M0[608], M0[579], M0[578], M0[31], M0[30]};
layer1_N21 layer1_N21_inst (.M0(layer1_N21_wire), .M1(M1[43:42]));

wire [11:0] layer1_N22_wire = {M0[615], M0[614], M0[529], M0[528], M0[523], M0[522], M0[453], M0[452], M0[383], M0[382], M0[271], M0[270]};
layer1_N22 layer1_N22_inst (.M0(layer1_N22_wire), .M1(M1[45:44]));

wire [11:0] layer1_N23_wire = {M0[855], M0[854], M0[777], M0[776], M0[433], M0[432], M0[387], M0[386], M0[181], M0[180], M0[77], M0[76]};
layer1_N23 layer1_N23_inst (.M0(layer1_N23_wire), .M1(M1[47:46]));

wire [11:0] layer1_N24_wire = {M0[1005], M0[1004], M0[945], M0[944], M0[861], M0[860], M0[547], M0[546], M0[413], M0[412], M0[29], M0[28]};
layer1_N24 layer1_N24_inst (.M0(layer1_N24_wire), .M1(M1[49:48]));

wire [11:0] layer1_N25_wire = {M0[749], M0[748], M0[619], M0[618], M0[435], M0[434], M0[429], M0[428], M0[53], M0[52], M0[11], M0[10]};
layer1_N25 layer1_N25_inst (.M0(layer1_N25_wire), .M1(M1[51:50]));

wire [11:0] layer1_N26_wire = {M0[1007], M0[1006], M0[559], M0[558], M0[341], M0[340], M0[241], M0[240], M0[21], M0[20], M0[5], M0[4]};
layer1_N26 layer1_N26_inst (.M0(layer1_N26_wire), .M1(M1[53:52]));

wire [11:0] layer1_N27_wire = {M0[843], M0[842], M0[659], M0[658], M0[485], M0[484], M0[171], M0[170], M0[119], M0[118], M0[23], M0[22]};
layer1_N27 layer1_N27_inst (.M0(layer1_N27_wire), .M1(M1[55:54]));

wire [11:0] layer1_N28_wire = {M0[997], M0[996], M0[791], M0[790], M0[407], M0[406], M0[353], M0[352], M0[115], M0[114], M0[111], M0[110]};
layer1_N28 layer1_N28_inst (.M0(layer1_N28_wire), .M1(M1[57:56]));

wire [11:0] layer1_N29_wire = {M0[895], M0[894], M0[835], M0[834], M0[623], M0[622], M0[269], M0[268], M0[253], M0[252], M0[149], M0[148]};
layer1_N29 layer1_N29_inst (.M0(layer1_N29_wire), .M1(M1[59:58]));

wire [11:0] layer1_N30_wire = {M0[597], M0[596], M0[571], M0[570], M0[483], M0[482], M0[385], M0[384], M0[203], M0[202], M0[199], M0[198]};
layer1_N30 layer1_N30_inst (.M0(layer1_N30_wire), .M1(M1[61:60]));

wire [11:0] layer1_N31_wire = {M0[767], M0[766], M0[729], M0[728], M0[503], M0[502], M0[269], M0[268], M0[203], M0[202], M0[91], M0[90]};
layer1_N31 layer1_N31_inst (.M0(layer1_N31_wire), .M1(M1[63:62]));

wire [11:0] layer1_N32_wire = {M0[983], M0[982], M0[863], M0[862], M0[617], M0[616], M0[517], M0[516], M0[287], M0[286], M0[273], M0[272]};
layer1_N32 layer1_N32_inst (.M0(layer1_N32_wire), .M1(M1[65:64]));

wire [11:0] layer1_N33_wire = {M0[995], M0[994], M0[923], M0[922], M0[703], M0[702], M0[677], M0[676], M0[99], M0[98], M0[43], M0[42]};
layer1_N33 layer1_N33_inst (.M0(layer1_N33_wire), .M1(M1[67:66]));

wire [11:0] layer1_N34_wire = {M0[923], M0[922], M0[881], M0[880], M0[799], M0[798], M0[545], M0[544], M0[137], M0[136], M0[45], M0[44]};
layer1_N34 layer1_N34_inst (.M0(layer1_N34_wire), .M1(M1[69:68]));

wire [11:0] layer1_N35_wire = {M0[871], M0[870], M0[797], M0[796], M0[495], M0[494], M0[437], M0[436], M0[227], M0[226], M0[93], M0[92]};
layer1_N35 layer1_N35_inst (.M0(layer1_N35_wire), .M1(M1[71:70]));

wire [11:0] layer1_N36_wire = {M0[547], M0[546], M0[399], M0[398], M0[389], M0[388], M0[307], M0[306], M0[167], M0[166], M0[143], M0[142]};
layer1_N36 layer1_N36_inst (.M0(layer1_N36_wire), .M1(M1[73:72]));

wire [11:0] layer1_N37_wire = {M0[943], M0[942], M0[751], M0[750], M0[645], M0[644], M0[597], M0[596], M0[457], M0[456], M0[13], M0[12]};
layer1_N37 layer1_N37_inst (.M0(layer1_N37_wire), .M1(M1[75:74]));

wire [11:0] layer1_N38_wire = {M0[847], M0[846], M0[575], M0[574], M0[503], M0[502], M0[497], M0[496], M0[357], M0[356], M0[323], M0[322]};
layer1_N38 layer1_N38_inst (.M0(layer1_N38_wire), .M1(M1[77:76]));

wire [11:0] layer1_N39_wire = {M0[573], M0[572], M0[499], M0[498], M0[455], M0[454], M0[305], M0[304], M0[183], M0[182], M0[27], M0[26]};
layer1_N39 layer1_N39_inst (.M0(layer1_N39_wire), .M1(M1[79:78]));

wire [11:0] layer1_N40_wire = {M0[1007], M0[1006], M0[957], M0[956], M0[739], M0[738], M0[479], M0[478], M0[325], M0[324], M0[119], M0[118]};
layer1_N40 layer1_N40_inst (.M0(layer1_N40_wire), .M1(M1[81:80]));

wire [11:0] layer1_N41_wire = {M0[953], M0[952], M0[897], M0[896], M0[811], M0[810], M0[517], M0[516], M0[297], M0[296], M0[125], M0[124]};
layer1_N41 layer1_N41_inst (.M0(layer1_N41_wire), .M1(M1[83:82]));

wire [11:0] layer1_N42_wire = {M0[1005], M0[1004], M0[487], M0[486], M0[315], M0[314], M0[297], M0[296], M0[105], M0[104], M0[79], M0[78]};
layer1_N42 layer1_N42_inst (.M0(layer1_N42_wire), .M1(M1[85:84]));

wire [11:0] layer1_N43_wire = {M0[935], M0[934], M0[811], M0[810], M0[805], M0[804], M0[747], M0[746], M0[735], M0[734], M0[489], M0[488]};
layer1_N43 layer1_N43_inst (.M0(layer1_N43_wire), .M1(M1[87:86]));

wire [11:0] layer1_N44_wire = {M0[895], M0[894], M0[877], M0[876], M0[473], M0[472], M0[275], M0[274], M0[187], M0[186], M0[41], M0[40]};
layer1_N44 layer1_N44_inst (.M0(layer1_N44_wire), .M1(M1[89:88]));

wire [11:0] layer1_N45_wire = {M0[973], M0[972], M0[587], M0[586], M0[557], M0[556], M0[413], M0[412], M0[169], M0[168], M0[35], M0[34]};
layer1_N45 layer1_N45_inst (.M0(layer1_N45_wire), .M1(M1[91:90]));

wire [11:0] layer1_N46_wire = {M0[889], M0[888], M0[777], M0[776], M0[717], M0[716], M0[401], M0[400], M0[171], M0[170], M0[65], M0[64]};
layer1_N46 layer1_N46_inst (.M0(layer1_N46_wire), .M1(M1[93:92]));

wire [11:0] layer1_N47_wire = {M0[1021], M0[1020], M0[991], M0[990], M0[771], M0[770], M0[399], M0[398], M0[277], M0[276], M0[59], M0[58]};
layer1_N47 layer1_N47_inst (.M0(layer1_N47_wire), .M1(M1[95:94]));

wire [11:0] layer1_N48_wire = {M0[967], M0[966], M0[809], M0[808], M0[789], M0[788], M0[689], M0[688], M0[573], M0[572], M0[255], M0[254]};
layer1_N48 layer1_N48_inst (.M0(layer1_N48_wire), .M1(M1[97:96]));

wire [11:0] layer1_N49_wire = {M0[969], M0[968], M0[943], M0[942], M0[525], M0[524], M0[451], M0[450], M0[359], M0[358], M0[339], M0[338]};
layer1_N49 layer1_N49_inst (.M0(layer1_N49_wire), .M1(M1[99:98]));

wire [11:0] layer1_N50_wire = {M0[951], M0[950], M0[597], M0[596], M0[501], M0[500], M0[317], M0[316], M0[235], M0[234], M0[225], M0[224]};
layer1_N50 layer1_N50_inst (.M0(layer1_N50_wire), .M1(M1[101:100]));

wire [11:0] layer1_N51_wire = {M0[985], M0[984], M0[521], M0[520], M0[469], M0[468], M0[457], M0[456], M0[33], M0[32], M0[29], M0[28]};
layer1_N51 layer1_N51_inst (.M0(layer1_N51_wire), .M1(M1[103:102]));

wire [11:0] layer1_N52_wire = {M0[977], M0[976], M0[683], M0[682], M0[495], M0[494], M0[347], M0[346], M0[101], M0[100], M0[23], M0[22]};
layer1_N52 layer1_N52_inst (.M0(layer1_N52_wire), .M1(M1[105:104]));

wire [11:0] layer1_N53_wire = {M0[757], M0[756], M0[721], M0[720], M0[531], M0[530], M0[289], M0[288], M0[195], M0[194], M0[145], M0[144]};
layer1_N53 layer1_N53_inst (.M0(layer1_N53_wire), .M1(M1[107:106]));

wire [11:0] layer1_N54_wire = {M0[863], M0[862], M0[775], M0[774], M0[421], M0[420], M0[297], M0[296], M0[281], M0[280], M0[17], M0[16]};
layer1_N54 layer1_N54_inst (.M0(layer1_N54_wire), .M1(M1[109:108]));

wire [11:0] layer1_N55_wire = {M0[987], M0[986], M0[459], M0[458], M0[401], M0[400], M0[141], M0[140], M0[95], M0[94], M0[19], M0[18]};
layer1_N55 layer1_N55_inst (.M0(layer1_N55_wire), .M1(M1[111:110]));

wire [11:0] layer1_N56_wire = {M0[915], M0[914], M0[837], M0[836], M0[345], M0[344], M0[309], M0[308], M0[97], M0[96], M0[65], M0[64]};
layer1_N56 layer1_N56_inst (.M0(layer1_N56_wire), .M1(M1[113:112]));

wire [11:0] layer1_N57_wire = {M0[799], M0[798], M0[759], M0[758], M0[613], M0[612], M0[567], M0[566], M0[529], M0[528], M0[287], M0[286]};
layer1_N57 layer1_N57_inst (.M0(layer1_N57_wire), .M1(M1[115:114]));

wire [11:0] layer1_N58_wire = {M0[725], M0[724], M0[683], M0[682], M0[341], M0[340], M0[319], M0[318], M0[193], M0[192], M0[153], M0[152]};
layer1_N58 layer1_N58_inst (.M0(layer1_N58_wire), .M1(M1[117:116]));

wire [11:0] layer1_N59_wire = {M0[855], M0[854], M0[775], M0[774], M0[713], M0[712], M0[317], M0[316], M0[243], M0[242], M0[81], M0[80]};
layer1_N59 layer1_N59_inst (.M0(layer1_N59_wire), .M1(M1[119:118]));

wire [11:0] layer1_N60_wire = {M0[907], M0[906], M0[315], M0[314], M0[127], M0[126], M0[99], M0[98], M0[91], M0[90], M0[81], M0[80]};
layer1_N60 layer1_N60_inst (.M0(layer1_N60_wire), .M1(M1[121:120]));

wire [11:0] layer1_N61_wire = {M0[1023], M0[1022], M0[827], M0[826], M0[535], M0[534], M0[195], M0[194], M0[115], M0[114], M0[73], M0[72]};
layer1_N61 layer1_N61_inst (.M0(layer1_N61_wire), .M1(M1[123:122]));

wire [11:0] layer1_N62_wire = {M0[647], M0[646], M0[611], M0[610], M0[585], M0[584], M0[523], M0[522], M0[471], M0[470], M0[291], M0[290]};
layer1_N62 layer1_N62_inst (.M0(layer1_N62_wire), .M1(M1[125:124]));

wire [11:0] layer1_N63_wire = {M0[887], M0[886], M0[795], M0[794], M0[765], M0[764], M0[693], M0[692], M0[529], M0[528], M0[507], M0[506]};
layer1_N63 layer1_N63_inst (.M0(layer1_N63_wire), .M1(M1[127:126]));

wire [11:0] layer1_N64_wire = {M0[763], M0[762], M0[561], M0[560], M0[539], M0[538], M0[363], M0[362], M0[37], M0[36], M0[23], M0[22]};
layer1_N64 layer1_N64_inst (.M0(layer1_N64_wire), .M1(M1[129:128]));

wire [11:0] layer1_N65_wire = {M0[639], M0[638], M0[625], M0[624], M0[261], M0[260], M0[241], M0[240], M0[205], M0[204], M0[17], M0[16]};
layer1_N65 layer1_N65_inst (.M0(layer1_N65_wire), .M1(M1[131:130]));

wire [11:0] layer1_N66_wire = {M0[789], M0[788], M0[693], M0[692], M0[635], M0[634], M0[523], M0[522], M0[395], M0[394], M0[25], M0[24]};
layer1_N66 layer1_N66_inst (.M0(layer1_N66_wire), .M1(M1[133:132]));

wire [11:0] layer1_N67_wire = {M0[807], M0[806], M0[781], M0[780], M0[675], M0[674], M0[625], M0[624], M0[505], M0[504], M0[489], M0[488]};
layer1_N67 layer1_N67_inst (.M0(layer1_N67_wire), .M1(M1[135:134]));

wire [11:0] layer1_N68_wire = {M0[1009], M0[1008], M0[739], M0[738], M0[727], M0[726], M0[301], M0[300], M0[233], M0[232], M0[149], M0[148]};
layer1_N68 layer1_N68_inst (.M0(layer1_N68_wire), .M1(M1[137:136]));

wire [11:0] layer1_N69_wire = {M0[997], M0[996], M0[927], M0[926], M0[845], M0[844], M0[711], M0[710], M0[523], M0[522], M0[139], M0[138]};
layer1_N69 layer1_N69_inst (.M0(layer1_N69_wire), .M1(M1[139:138]));

wire [11:0] layer1_N70_wire = {M0[887], M0[886], M0[743], M0[742], M0[493], M0[492], M0[485], M0[484], M0[387], M0[386], M0[375], M0[374]};
layer1_N70 layer1_N70_inst (.M0(layer1_N70_wire), .M1(M1[141:140]));

wire [11:0] layer1_N71_wire = {M0[839], M0[838], M0[773], M0[772], M0[765], M0[764], M0[725], M0[724], M0[383], M0[382], M0[45], M0[44]};
layer1_N71 layer1_N71_inst (.M0(layer1_N71_wire), .M1(M1[143:142]));

wire [11:0] layer1_N72_wire = {M0[967], M0[966], M0[875], M0[874], M0[867], M0[866], M0[751], M0[750], M0[271], M0[270], M0[65], M0[64]};
layer1_N72 layer1_N72_inst (.M0(layer1_N72_wire), .M1(M1[145:144]));

wire [11:0] layer1_N73_wire = {M0[945], M0[944], M0[825], M0[824], M0[777], M0[776], M0[273], M0[272], M0[175], M0[174], M0[141], M0[140]};
layer1_N73 layer1_N73_inst (.M0(layer1_N73_wire), .M1(M1[147:146]));

wire [11:0] layer1_N74_wire = {M0[609], M0[608], M0[479], M0[478], M0[187], M0[186], M0[175], M0[174], M0[123], M0[122], M0[37], M0[36]};
layer1_N74 layer1_N74_inst (.M0(layer1_N74_wire), .M1(M1[149:148]));

wire [11:0] layer1_N75_wire = {M0[867], M0[866], M0[715], M0[714], M0[473], M0[472], M0[331], M0[330], M0[193], M0[192], M0[73], M0[72]};
layer1_N75 layer1_N75_inst (.M0(layer1_N75_wire), .M1(M1[151:150]));

wire [11:0] layer1_N76_wire = {M0[761], M0[760], M0[643], M0[642], M0[285], M0[284], M0[165], M0[164], M0[39], M0[38], M0[25], M0[24]};
layer1_N76 layer1_N76_inst (.M0(layer1_N76_wire), .M1(M1[153:152]));

wire [11:0] layer1_N77_wire = {M0[875], M0[874], M0[669], M0[668], M0[559], M0[558], M0[379], M0[378], M0[117], M0[116], M0[51], M0[50]};
layer1_N77 layer1_N77_inst (.M0(layer1_N77_wire), .M1(M1[155:154]));

wire [11:0] layer1_N78_wire = {M0[935], M0[934], M0[753], M0[752], M0[713], M0[712], M0[677], M0[676], M0[239], M0[238], M0[183], M0[182]};
layer1_N78 layer1_N78_inst (.M0(layer1_N78_wire), .M1(M1[157:156]));

wire [11:0] layer1_N79_wire = {M0[679], M0[678], M0[631], M0[630], M0[425], M0[424], M0[299], M0[298], M0[249], M0[248], M0[71], M0[70]};
layer1_N79 layer1_N79_inst (.M0(layer1_N79_wire), .M1(M1[159:158]));

wire [11:0] layer1_N80_wire = {M0[433], M0[432], M0[303], M0[302], M0[213], M0[212], M0[123], M0[122], M0[69], M0[68], M0[29], M0[28]};
layer1_N80 layer1_N80_inst (.M0(layer1_N80_wire), .M1(M1[161:160]));

wire [11:0] layer1_N81_wire = {M0[1023], M0[1022], M0[783], M0[782], M0[473], M0[472], M0[295], M0[294], M0[151], M0[150], M0[55], M0[54]};
layer1_N81 layer1_N81_inst (.M0(layer1_N81_wire), .M1(M1[163:162]));

wire [11:0] layer1_N82_wire = {M0[853], M0[852], M0[691], M0[690], M0[377], M0[376], M0[309], M0[308], M0[219], M0[218], M0[3], M0[2]};
layer1_N82 layer1_N82_inst (.M0(layer1_N82_wire), .M1(M1[165:164]));

wire [11:0] layer1_N83_wire = {M0[959], M0[958], M0[861], M0[860], M0[769], M0[768], M0[631], M0[630], M0[557], M0[556], M0[501], M0[500]};
layer1_N83 layer1_N83_inst (.M0(layer1_N83_wire), .M1(M1[167:166]));

wire [11:0] layer1_N84_wire = {M0[953], M0[952], M0[739], M0[738], M0[707], M0[706], M0[479], M0[478], M0[355], M0[354], M0[77], M0[76]};
layer1_N84 layer1_N84_inst (.M0(layer1_N84_wire), .M1(M1[169:168]));

wire [11:0] layer1_N85_wire = {M0[877], M0[876], M0[777], M0[776], M0[755], M0[754], M0[491], M0[490], M0[21], M0[20], M0[3], M0[2]};
layer1_N85 layer1_N85_inst (.M0(layer1_N85_wire), .M1(M1[171:170]));

endmodule