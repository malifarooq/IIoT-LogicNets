module layer3_N5 ( input [13:0] M0, output [1:0] M1 );

	(*rom_style = "distributed" *) reg [1:0] M1r;
	assign M1 = M1r;
	always @ (M0) begin
		case (M0)
			14'b00000000000000: M1r = 2'b00;
			14'b01000000000000: M1r = 2'b00;
			14'b10000000000000: M1r = 2'b00;
			14'b11000000000000: M1r = 2'b00;
			14'b00010000000000: M1r = 2'b00;
			14'b01010000000000: M1r = 2'b00;
			14'b10010000000000: M1r = 2'b00;
			14'b11010000000000: M1r = 2'b00;
			14'b00100000000000: M1r = 2'b00;
			14'b01100000000000: M1r = 2'b00;
			14'b10100000000000: M1r = 2'b00;
			14'b11100000000000: M1r = 2'b00;
			14'b00110000000000: M1r = 2'b00;
			14'b01110000000000: M1r = 2'b00;
			14'b10110000000000: M1r = 2'b00;
			14'b11110000000000: M1r = 2'b00;
			14'b00000100000000: M1r = 2'b00;
			14'b01000100000000: M1r = 2'b00;
			14'b10000100000000: M1r = 2'b00;
			14'b11000100000000: M1r = 2'b00;
			14'b00010100000000: M1r = 2'b00;
			14'b01010100000000: M1r = 2'b00;
			14'b10010100000000: M1r = 2'b00;
			14'b11010100000000: M1r = 2'b00;
			14'b00100100000000: M1r = 2'b00;
			14'b01100100000000: M1r = 2'b00;
			14'b10100100000000: M1r = 2'b00;
			14'b11100100000000: M1r = 2'b00;
			14'b00110100000000: M1r = 2'b00;
			14'b01110100000000: M1r = 2'b00;
			14'b10110100000000: M1r = 2'b00;
			14'b11110100000000: M1r = 2'b00;
			14'b00001000000000: M1r = 2'b01;
			14'b01001000000000: M1r = 2'b01;
			14'b10001000000000: M1r = 2'b01;
			14'b11001000000000: M1r = 2'b01;
			14'b00011000000000: M1r = 2'b00;
			14'b01011000000000: M1r = 2'b00;
			14'b10011000000000: M1r = 2'b00;
			14'b11011000000000: M1r = 2'b01;
			14'b00101000000000: M1r = 2'b00;
			14'b01101000000000: M1r = 2'b00;
			14'b10101000000000: M1r = 2'b00;
			14'b11101000000000: M1r = 2'b00;
			14'b00111000000000: M1r = 2'b00;
			14'b01111000000000: M1r = 2'b00;
			14'b10111000000000: M1r = 2'b00;
			14'b11111000000000: M1r = 2'b00;
			14'b00001100000000: M1r = 2'b01;
			14'b01001100000000: M1r = 2'b10;
			14'b10001100000000: M1r = 2'b10;
			14'b11001100000000: M1r = 2'b10;
			14'b00011100000000: M1r = 2'b01;
			14'b01011100000000: M1r = 2'b01;
			14'b10011100000000: M1r = 2'b01;
			14'b11011100000000: M1r = 2'b01;
			14'b00101100000000: M1r = 2'b00;
			14'b01101100000000: M1r = 2'b01;
			14'b10101100000000: M1r = 2'b01;
			14'b11101100000000: M1r = 2'b01;
			14'b00111100000000: M1r = 2'b00;
			14'b01111100000000: M1r = 2'b00;
			14'b10111100000000: M1r = 2'b00;
			14'b11111100000000: M1r = 2'b00;
			14'b00000001000000: M1r = 2'b00;
			14'b01000001000000: M1r = 2'b00;
			14'b10000001000000: M1r = 2'b00;
			14'b11000001000000: M1r = 2'b00;
			14'b00010001000000: M1r = 2'b00;
			14'b01010001000000: M1r = 2'b00;
			14'b10010001000000: M1r = 2'b00;
			14'b11010001000000: M1r = 2'b00;
			14'b00100001000000: M1r = 2'b00;
			14'b01100001000000: M1r = 2'b00;
			14'b10100001000000: M1r = 2'b00;
			14'b11100001000000: M1r = 2'b00;
			14'b00110001000000: M1r = 2'b00;
			14'b01110001000000: M1r = 2'b00;
			14'b10110001000000: M1r = 2'b00;
			14'b11110001000000: M1r = 2'b00;
			14'b00000101000000: M1r = 2'b00;
			14'b01000101000000: M1r = 2'b00;
			14'b10000101000000: M1r = 2'b00;
			14'b11000101000000: M1r = 2'b00;
			14'b00010101000000: M1r = 2'b00;
			14'b01010101000000: M1r = 2'b00;
			14'b10010101000000: M1r = 2'b00;
			14'b11010101000000: M1r = 2'b00;
			14'b00100101000000: M1r = 2'b00;
			14'b01100101000000: M1r = 2'b00;
			14'b10100101000000: M1r = 2'b00;
			14'b11100101000000: M1r = 2'b00;
			14'b00110101000000: M1r = 2'b00;
			14'b01110101000000: M1r = 2'b00;
			14'b10110101000000: M1r = 2'b00;
			14'b11110101000000: M1r = 2'b00;
			14'b00001001000000: M1r = 2'b00;
			14'b01001001000000: M1r = 2'b01;
			14'b10001001000000: M1r = 2'b01;
			14'b11001001000000: M1r = 2'b01;
			14'b00011001000000: M1r = 2'b00;
			14'b01011001000000: M1r = 2'b00;
			14'b10011001000000: M1r = 2'b00;
			14'b11011001000000: M1r = 2'b00;
			14'b00101001000000: M1r = 2'b00;
			14'b01101001000000: M1r = 2'b00;
			14'b10101001000000: M1r = 2'b00;
			14'b11101001000000: M1r = 2'b00;
			14'b00111001000000: M1r = 2'b00;
			14'b01111001000000: M1r = 2'b00;
			14'b10111001000000: M1r = 2'b00;
			14'b11111001000000: M1r = 2'b00;
			14'b00001101000000: M1r = 2'b01;
			14'b01001101000000: M1r = 2'b01;
			14'b10001101000000: M1r = 2'b01;
			14'b11001101000000: M1r = 2'b10;
			14'b00011101000000: M1r = 2'b01;
			14'b01011101000000: M1r = 2'b01;
			14'b10011101000000: M1r = 2'b01;
			14'b11011101000000: M1r = 2'b01;
			14'b00101101000000: M1r = 2'b00;
			14'b01101101000000: M1r = 2'b00;
			14'b10101101000000: M1r = 2'b00;
			14'b11101101000000: M1r = 2'b01;
			14'b00111101000000: M1r = 2'b00;
			14'b01111101000000: M1r = 2'b00;
			14'b10111101000000: M1r = 2'b00;
			14'b11111101000000: M1r = 2'b00;
			14'b00000010000000: M1r = 2'b00;
			14'b01000010000000: M1r = 2'b00;
			14'b10000010000000: M1r = 2'b00;
			14'b11000010000000: M1r = 2'b00;
			14'b00010010000000: M1r = 2'b00;
			14'b01010010000000: M1r = 2'b00;
			14'b10010010000000: M1r = 2'b00;
			14'b11010010000000: M1r = 2'b00;
			14'b00100010000000: M1r = 2'b00;
			14'b01100010000000: M1r = 2'b00;
			14'b10100010000000: M1r = 2'b00;
			14'b11100010000000: M1r = 2'b00;
			14'b00110010000000: M1r = 2'b00;
			14'b01110010000000: M1r = 2'b00;
			14'b10110010000000: M1r = 2'b00;
			14'b11110010000000: M1r = 2'b00;
			14'b00000110000000: M1r = 2'b00;
			14'b01000110000000: M1r = 2'b00;
			14'b10000110000000: M1r = 2'b00;
			14'b11000110000000: M1r = 2'b00;
			14'b00010110000000: M1r = 2'b00;
			14'b01010110000000: M1r = 2'b00;
			14'b10010110000000: M1r = 2'b00;
			14'b11010110000000: M1r = 2'b00;
			14'b00100110000000: M1r = 2'b00;
			14'b01100110000000: M1r = 2'b00;
			14'b10100110000000: M1r = 2'b00;
			14'b11100110000000: M1r = 2'b00;
			14'b00110110000000: M1r = 2'b00;
			14'b01110110000000: M1r = 2'b00;
			14'b10110110000000: M1r = 2'b00;
			14'b11110110000000: M1r = 2'b00;
			14'b00001010000000: M1r = 2'b00;
			14'b01001010000000: M1r = 2'b00;
			14'b10001010000000: M1r = 2'b00;
			14'b11001010000000: M1r = 2'b01;
			14'b00011010000000: M1r = 2'b00;
			14'b01011010000000: M1r = 2'b00;
			14'b10011010000000: M1r = 2'b00;
			14'b11011010000000: M1r = 2'b00;
			14'b00101010000000: M1r = 2'b00;
			14'b01101010000000: M1r = 2'b00;
			14'b10101010000000: M1r = 2'b00;
			14'b11101010000000: M1r = 2'b00;
			14'b00111010000000: M1r = 2'b00;
			14'b01111010000000: M1r = 2'b00;
			14'b10111010000000: M1r = 2'b00;
			14'b11111010000000: M1r = 2'b00;
			14'b00001110000000: M1r = 2'b01;
			14'b01001110000000: M1r = 2'b01;
			14'b10001110000000: M1r = 2'b01;
			14'b11001110000000: M1r = 2'b01;
			14'b00011110000000: M1r = 2'b00;
			14'b01011110000000: M1r = 2'b01;
			14'b10011110000000: M1r = 2'b01;
			14'b11011110000000: M1r = 2'b01;
			14'b00101110000000: M1r = 2'b00;
			14'b01101110000000: M1r = 2'b00;
			14'b10101110000000: M1r = 2'b00;
			14'b11101110000000: M1r = 2'b00;
			14'b00111110000000: M1r = 2'b00;
			14'b01111110000000: M1r = 2'b00;
			14'b10111110000000: M1r = 2'b00;
			14'b11111110000000: M1r = 2'b00;
			14'b00000011000000: M1r = 2'b00;
			14'b01000011000000: M1r = 2'b00;
			14'b10000011000000: M1r = 2'b00;
			14'b11000011000000: M1r = 2'b00;
			14'b00010011000000: M1r = 2'b00;
			14'b01010011000000: M1r = 2'b00;
			14'b10010011000000: M1r = 2'b00;
			14'b11010011000000: M1r = 2'b00;
			14'b00100011000000: M1r = 2'b00;
			14'b01100011000000: M1r = 2'b00;
			14'b10100011000000: M1r = 2'b00;
			14'b11100011000000: M1r = 2'b00;
			14'b00110011000000: M1r = 2'b00;
			14'b01110011000000: M1r = 2'b00;
			14'b10110011000000: M1r = 2'b00;
			14'b11110011000000: M1r = 2'b00;
			14'b00000111000000: M1r = 2'b00;
			14'b01000111000000: M1r = 2'b00;
			14'b10000111000000: M1r = 2'b00;
			14'b11000111000000: M1r = 2'b00;
			14'b00010111000000: M1r = 2'b00;
			14'b01010111000000: M1r = 2'b00;
			14'b10010111000000: M1r = 2'b00;
			14'b11010111000000: M1r = 2'b00;
			14'b00100111000000: M1r = 2'b00;
			14'b01100111000000: M1r = 2'b00;
			14'b10100111000000: M1r = 2'b00;
			14'b11100111000000: M1r = 2'b00;
			14'b00110111000000: M1r = 2'b00;
			14'b01110111000000: M1r = 2'b00;
			14'b10110111000000: M1r = 2'b00;
			14'b11110111000000: M1r = 2'b00;
			14'b00001011000000: M1r = 2'b00;
			14'b01001011000000: M1r = 2'b00;
			14'b10001011000000: M1r = 2'b00;
			14'b11001011000000: M1r = 2'b00;
			14'b00011011000000: M1r = 2'b00;
			14'b01011011000000: M1r = 2'b00;
			14'b10011011000000: M1r = 2'b00;
			14'b11011011000000: M1r = 2'b00;
			14'b00101011000000: M1r = 2'b00;
			14'b01101011000000: M1r = 2'b00;
			14'b10101011000000: M1r = 2'b00;
			14'b11101011000000: M1r = 2'b00;
			14'b00111011000000: M1r = 2'b00;
			14'b01111011000000: M1r = 2'b00;
			14'b10111011000000: M1r = 2'b00;
			14'b11111011000000: M1r = 2'b00;
			14'b00001111000000: M1r = 2'b01;
			14'b01001111000000: M1r = 2'b01;
			14'b10001111000000: M1r = 2'b01;
			14'b11001111000000: M1r = 2'b01;
			14'b00011111000000: M1r = 2'b00;
			14'b01011111000000: M1r = 2'b00;
			14'b10011111000000: M1r = 2'b00;
			14'b11011111000000: M1r = 2'b01;
			14'b00101111000000: M1r = 2'b00;
			14'b01101111000000: M1r = 2'b00;
			14'b10101111000000: M1r = 2'b00;
			14'b11101111000000: M1r = 2'b00;
			14'b00111111000000: M1r = 2'b00;
			14'b01111111000000: M1r = 2'b00;
			14'b10111111000000: M1r = 2'b00;
			14'b11111111000000: M1r = 2'b00;
			14'b00000000010000: M1r = 2'b00;
			14'b01000000010000: M1r = 2'b00;
			14'b10000000010000: M1r = 2'b00;
			14'b11000000010000: M1r = 2'b00;
			14'b00010000010000: M1r = 2'b00;
			14'b01010000010000: M1r = 2'b00;
			14'b10010000010000: M1r = 2'b00;
			14'b11010000010000: M1r = 2'b00;
			14'b00100000010000: M1r = 2'b00;
			14'b01100000010000: M1r = 2'b00;
			14'b10100000010000: M1r = 2'b00;
			14'b11100000010000: M1r = 2'b00;
			14'b00110000010000: M1r = 2'b00;
			14'b01110000010000: M1r = 2'b00;
			14'b10110000010000: M1r = 2'b00;
			14'b11110000010000: M1r = 2'b00;
			14'b00000100010000: M1r = 2'b00;
			14'b01000100010000: M1r = 2'b00;
			14'b10000100010000: M1r = 2'b01;
			14'b11000100010000: M1r = 2'b01;
			14'b00010100010000: M1r = 2'b00;
			14'b01010100010000: M1r = 2'b00;
			14'b10010100010000: M1r = 2'b00;
			14'b11010100010000: M1r = 2'b00;
			14'b00100100010000: M1r = 2'b00;
			14'b01100100010000: M1r = 2'b00;
			14'b10100100010000: M1r = 2'b00;
			14'b11100100010000: M1r = 2'b00;
			14'b00110100010000: M1r = 2'b00;
			14'b01110100010000: M1r = 2'b00;
			14'b10110100010000: M1r = 2'b00;
			14'b11110100010000: M1r = 2'b00;
			14'b00001000010000: M1r = 2'b01;
			14'b01001000010000: M1r = 2'b01;
			14'b10001000010000: M1r = 2'b01;
			14'b11001000010000: M1r = 2'b10;
			14'b00011000010000: M1r = 2'b01;
			14'b01011000010000: M1r = 2'b01;
			14'b10011000010000: M1r = 2'b01;
			14'b11011000010000: M1r = 2'b01;
			14'b00101000010000: M1r = 2'b00;
			14'b01101000010000: M1r = 2'b00;
			14'b10101000010000: M1r = 2'b00;
			14'b11101000010000: M1r = 2'b01;
			14'b00111000010000: M1r = 2'b00;
			14'b01111000010000: M1r = 2'b00;
			14'b10111000010000: M1r = 2'b00;
			14'b11111000010000: M1r = 2'b00;
			14'b00001100010000: M1r = 2'b10;
			14'b01001100010000: M1r = 2'b10;
			14'b10001100010000: M1r = 2'b10;
			14'b11001100010000: M1r = 2'b10;
			14'b00011100010000: M1r = 2'b01;
			14'b01011100010000: M1r = 2'b01;
			14'b10011100010000: M1r = 2'b10;
			14'b11011100010000: M1r = 2'b10;
			14'b00101100010000: M1r = 2'b01;
			14'b01101100010000: M1r = 2'b01;
			14'b10101100010000: M1r = 2'b01;
			14'b11101100010000: M1r = 2'b01;
			14'b00111100010000: M1r = 2'b00;
			14'b01111100010000: M1r = 2'b01;
			14'b10111100010000: M1r = 2'b01;
			14'b11111100010000: M1r = 2'b01;
			14'b00000001010000: M1r = 2'b00;
			14'b01000001010000: M1r = 2'b00;
			14'b10000001010000: M1r = 2'b00;
			14'b11000001010000: M1r = 2'b00;
			14'b00010001010000: M1r = 2'b00;
			14'b01010001010000: M1r = 2'b00;
			14'b10010001010000: M1r = 2'b00;
			14'b11010001010000: M1r = 2'b00;
			14'b00100001010000: M1r = 2'b00;
			14'b01100001010000: M1r = 2'b00;
			14'b10100001010000: M1r = 2'b00;
			14'b11100001010000: M1r = 2'b00;
			14'b00110001010000: M1r = 2'b00;
			14'b01110001010000: M1r = 2'b00;
			14'b10110001010000: M1r = 2'b00;
			14'b11110001010000: M1r = 2'b00;
			14'b00000101010000: M1r = 2'b00;
			14'b01000101010000: M1r = 2'b00;
			14'b10000101010000: M1r = 2'b00;
			14'b11000101010000: M1r = 2'b01;
			14'b00010101010000: M1r = 2'b00;
			14'b01010101010000: M1r = 2'b00;
			14'b10010101010000: M1r = 2'b00;
			14'b11010101010000: M1r = 2'b00;
			14'b00100101010000: M1r = 2'b00;
			14'b01100101010000: M1r = 2'b00;
			14'b10100101010000: M1r = 2'b00;
			14'b11100101010000: M1r = 2'b00;
			14'b00110101010000: M1r = 2'b00;
			14'b01110101010000: M1r = 2'b00;
			14'b10110101010000: M1r = 2'b00;
			14'b11110101010000: M1r = 2'b00;
			14'b00001001010000: M1r = 2'b01;
			14'b01001001010000: M1r = 2'b01;
			14'b10001001010000: M1r = 2'b01;
			14'b11001001010000: M1r = 2'b01;
			14'b00011001010000: M1r = 2'b00;
			14'b01011001010000: M1r = 2'b00;
			14'b10011001010000: M1r = 2'b01;
			14'b11011001010000: M1r = 2'b01;
			14'b00101001010000: M1r = 2'b00;
			14'b01101001010000: M1r = 2'b00;
			14'b10101001010000: M1r = 2'b00;
			14'b11101001010000: M1r = 2'b00;
			14'b00111001010000: M1r = 2'b00;
			14'b01111001010000: M1r = 2'b00;
			14'b10111001010000: M1r = 2'b00;
			14'b11111001010000: M1r = 2'b00;
			14'b00001101010000: M1r = 2'b10;
			14'b01001101010000: M1r = 2'b10;
			14'b10001101010000: M1r = 2'b10;
			14'b11001101010000: M1r = 2'b10;
			14'b00011101010000: M1r = 2'b01;
			14'b01011101010000: M1r = 2'b01;
			14'b10011101010000: M1r = 2'b01;
			14'b11011101010000: M1r = 2'b10;
			14'b00101101010000: M1r = 2'b01;
			14'b01101101010000: M1r = 2'b01;
			14'b10101101010000: M1r = 2'b01;
			14'b11101101010000: M1r = 2'b01;
			14'b00111101010000: M1r = 2'b00;
			14'b01111101010000: M1r = 2'b00;
			14'b10111101010000: M1r = 2'b00;
			14'b11111101010000: M1r = 2'b01;
			14'b00000010010000: M1r = 2'b00;
			14'b01000010010000: M1r = 2'b00;
			14'b10000010010000: M1r = 2'b00;
			14'b11000010010000: M1r = 2'b00;
			14'b00010010010000: M1r = 2'b00;
			14'b01010010010000: M1r = 2'b00;
			14'b10010010010000: M1r = 2'b00;
			14'b11010010010000: M1r = 2'b00;
			14'b00100010010000: M1r = 2'b00;
			14'b01100010010000: M1r = 2'b00;
			14'b10100010010000: M1r = 2'b00;
			14'b11100010010000: M1r = 2'b00;
			14'b00110010010000: M1r = 2'b00;
			14'b01110010010000: M1r = 2'b00;
			14'b10110010010000: M1r = 2'b00;
			14'b11110010010000: M1r = 2'b00;
			14'b00000110010000: M1r = 2'b00;
			14'b01000110010000: M1r = 2'b00;
			14'b10000110010000: M1r = 2'b00;
			14'b11000110010000: M1r = 2'b00;
			14'b00010110010000: M1r = 2'b00;
			14'b01010110010000: M1r = 2'b00;
			14'b10010110010000: M1r = 2'b00;
			14'b11010110010000: M1r = 2'b00;
			14'b00100110010000: M1r = 2'b00;
			14'b01100110010000: M1r = 2'b00;
			14'b10100110010000: M1r = 2'b00;
			14'b11100110010000: M1r = 2'b00;
			14'b00110110010000: M1r = 2'b00;
			14'b01110110010000: M1r = 2'b00;
			14'b10110110010000: M1r = 2'b00;
			14'b11110110010000: M1r = 2'b00;
			14'b00001010010000: M1r = 2'b01;
			14'b01001010010000: M1r = 2'b01;
			14'b10001010010000: M1r = 2'b01;
			14'b11001010010000: M1r = 2'b01;
			14'b00011010010000: M1r = 2'b00;
			14'b01011010010000: M1r = 2'b00;
			14'b10011010010000: M1r = 2'b00;
			14'b11011010010000: M1r = 2'b01;
			14'b00101010010000: M1r = 2'b00;
			14'b01101010010000: M1r = 2'b00;
			14'b10101010010000: M1r = 2'b00;
			14'b11101010010000: M1r = 2'b00;
			14'b00111010010000: M1r = 2'b00;
			14'b01111010010000: M1r = 2'b00;
			14'b10111010010000: M1r = 2'b00;
			14'b11111010010000: M1r = 2'b00;
			14'b00001110010000: M1r = 2'b01;
			14'b01001110010000: M1r = 2'b01;
			14'b10001110010000: M1r = 2'b10;
			14'b11001110010000: M1r = 2'b10;
			14'b00011110010000: M1r = 2'b01;
			14'b01011110010000: M1r = 2'b01;
			14'b10011110010000: M1r = 2'b01;
			14'b11011110010000: M1r = 2'b01;
			14'b00101110010000: M1r = 2'b00;
			14'b01101110010000: M1r = 2'b00;
			14'b10101110010000: M1r = 2'b01;
			14'b11101110010000: M1r = 2'b01;
			14'b00111110010000: M1r = 2'b00;
			14'b01111110010000: M1r = 2'b00;
			14'b10111110010000: M1r = 2'b00;
			14'b11111110010000: M1r = 2'b00;
			14'b00000011010000: M1r = 2'b00;
			14'b01000011010000: M1r = 2'b00;
			14'b10000011010000: M1r = 2'b00;
			14'b11000011010000: M1r = 2'b00;
			14'b00010011010000: M1r = 2'b00;
			14'b01010011010000: M1r = 2'b00;
			14'b10010011010000: M1r = 2'b00;
			14'b11010011010000: M1r = 2'b00;
			14'b00100011010000: M1r = 2'b00;
			14'b01100011010000: M1r = 2'b00;
			14'b10100011010000: M1r = 2'b00;
			14'b11100011010000: M1r = 2'b00;
			14'b00110011010000: M1r = 2'b00;
			14'b01110011010000: M1r = 2'b00;
			14'b10110011010000: M1r = 2'b00;
			14'b11110011010000: M1r = 2'b00;
			14'b00000111010000: M1r = 2'b00;
			14'b01000111010000: M1r = 2'b00;
			14'b10000111010000: M1r = 2'b00;
			14'b11000111010000: M1r = 2'b00;
			14'b00010111010000: M1r = 2'b00;
			14'b01010111010000: M1r = 2'b00;
			14'b10010111010000: M1r = 2'b00;
			14'b11010111010000: M1r = 2'b00;
			14'b00100111010000: M1r = 2'b00;
			14'b01100111010000: M1r = 2'b00;
			14'b10100111010000: M1r = 2'b00;
			14'b11100111010000: M1r = 2'b00;
			14'b00110111010000: M1r = 2'b00;
			14'b01110111010000: M1r = 2'b00;
			14'b10110111010000: M1r = 2'b00;
			14'b11110111010000: M1r = 2'b00;
			14'b00001011010000: M1r = 2'b00;
			14'b01001011010000: M1r = 2'b00;
			14'b10001011010000: M1r = 2'b01;
			14'b11001011010000: M1r = 2'b01;
			14'b00011011010000: M1r = 2'b00;
			14'b01011011010000: M1r = 2'b00;
			14'b10011011010000: M1r = 2'b00;
			14'b11011011010000: M1r = 2'b00;
			14'b00101011010000: M1r = 2'b00;
			14'b01101011010000: M1r = 2'b00;
			14'b10101011010000: M1r = 2'b00;
			14'b11101011010000: M1r = 2'b00;
			14'b00111011010000: M1r = 2'b00;
			14'b01111011010000: M1r = 2'b00;
			14'b10111011010000: M1r = 2'b00;
			14'b11111011010000: M1r = 2'b00;
			14'b00001111010000: M1r = 2'b01;
			14'b01001111010000: M1r = 2'b01;
			14'b10001111010000: M1r = 2'b01;
			14'b11001111010000: M1r = 2'b01;
			14'b00011111010000: M1r = 2'b01;
			14'b01011111010000: M1r = 2'b01;
			14'b10011111010000: M1r = 2'b01;
			14'b11011111010000: M1r = 2'b01;
			14'b00101111010000: M1r = 2'b00;
			14'b01101111010000: M1r = 2'b00;
			14'b10101111010000: M1r = 2'b00;
			14'b11101111010000: M1r = 2'b01;
			14'b00111111010000: M1r = 2'b00;
			14'b01111111010000: M1r = 2'b00;
			14'b10111111010000: M1r = 2'b00;
			14'b11111111010000: M1r = 2'b00;
			14'b00000000100000: M1r = 2'b00;
			14'b01000000100000: M1r = 2'b00;
			14'b10000000100000: M1r = 2'b00;
			14'b11000000100000: M1r = 2'b00;
			14'b00010000100000: M1r = 2'b00;
			14'b01010000100000: M1r = 2'b00;
			14'b10010000100000: M1r = 2'b00;
			14'b11010000100000: M1r = 2'b00;
			14'b00100000100000: M1r = 2'b00;
			14'b01100000100000: M1r = 2'b00;
			14'b10100000100000: M1r = 2'b00;
			14'b11100000100000: M1r = 2'b00;
			14'b00110000100000: M1r = 2'b00;
			14'b01110000100000: M1r = 2'b00;
			14'b10110000100000: M1r = 2'b00;
			14'b11110000100000: M1r = 2'b00;
			14'b00000100100000: M1r = 2'b01;
			14'b01000100100000: M1r = 2'b01;
			14'b10000100100000: M1r = 2'b01;
			14'b11000100100000: M1r = 2'b01;
			14'b00010100100000: M1r = 2'b00;
			14'b01010100100000: M1r = 2'b00;
			14'b10010100100000: M1r = 2'b01;
			14'b11010100100000: M1r = 2'b01;
			14'b00100100100000: M1r = 2'b00;
			14'b01100100100000: M1r = 2'b00;
			14'b10100100100000: M1r = 2'b00;
			14'b11100100100000: M1r = 2'b00;
			14'b00110100100000: M1r = 2'b00;
			14'b01110100100000: M1r = 2'b00;
			14'b10110100100000: M1r = 2'b00;
			14'b11110100100000: M1r = 2'b00;
			14'b00001000100000: M1r = 2'b01;
			14'b01001000100000: M1r = 2'b10;
			14'b10001000100000: M1r = 2'b10;
			14'b11001000100000: M1r = 2'b10;
			14'b00011000100000: M1r = 2'b01;
			14'b01011000100000: M1r = 2'b01;
			14'b10011000100000: M1r = 2'b01;
			14'b11011000100000: M1r = 2'b01;
			14'b00101000100000: M1r = 2'b01;
			14'b01101000100000: M1r = 2'b01;
			14'b10101000100000: M1r = 2'b01;
			14'b11101000100000: M1r = 2'b01;
			14'b00111000100000: M1r = 2'b00;
			14'b01111000100000: M1r = 2'b00;
			14'b10111000100000: M1r = 2'b00;
			14'b11111000100000: M1r = 2'b01;
			14'b00001100100000: M1r = 2'b10;
			14'b01001100100000: M1r = 2'b10;
			14'b10001100100000: M1r = 2'b11;
			14'b11001100100000: M1r = 2'b11;
			14'b00011100100000: M1r = 2'b10;
			14'b01011100100000: M1r = 2'b10;
			14'b10011100100000: M1r = 2'b10;
			14'b11011100100000: M1r = 2'b10;
			14'b00101100100000: M1r = 2'b01;
			14'b01101100100000: M1r = 2'b01;
			14'b10101100100000: M1r = 2'b10;
			14'b11101100100000: M1r = 2'b10;
			14'b00111100100000: M1r = 2'b01;
			14'b01111100100000: M1r = 2'b01;
			14'b10111100100000: M1r = 2'b01;
			14'b11111100100000: M1r = 2'b01;
			14'b00000001100000: M1r = 2'b00;
			14'b01000001100000: M1r = 2'b00;
			14'b10000001100000: M1r = 2'b00;
			14'b11000001100000: M1r = 2'b00;
			14'b00010001100000: M1r = 2'b00;
			14'b01010001100000: M1r = 2'b00;
			14'b10010001100000: M1r = 2'b00;
			14'b11010001100000: M1r = 2'b00;
			14'b00100001100000: M1r = 2'b00;
			14'b01100001100000: M1r = 2'b00;
			14'b10100001100000: M1r = 2'b00;
			14'b11100001100000: M1r = 2'b00;
			14'b00110001100000: M1r = 2'b00;
			14'b01110001100000: M1r = 2'b00;
			14'b10110001100000: M1r = 2'b00;
			14'b11110001100000: M1r = 2'b00;
			14'b00000101100000: M1r = 2'b00;
			14'b01000101100000: M1r = 2'b01;
			14'b10000101100000: M1r = 2'b01;
			14'b11000101100000: M1r = 2'b01;
			14'b00010101100000: M1r = 2'b00;
			14'b01010101100000: M1r = 2'b00;
			14'b10010101100000: M1r = 2'b00;
			14'b11010101100000: M1r = 2'b00;
			14'b00100101100000: M1r = 2'b00;
			14'b01100101100000: M1r = 2'b00;
			14'b10100101100000: M1r = 2'b00;
			14'b11100101100000: M1r = 2'b00;
			14'b00110101100000: M1r = 2'b00;
			14'b01110101100000: M1r = 2'b00;
			14'b10110101100000: M1r = 2'b00;
			14'b11110101100000: M1r = 2'b00;
			14'b00001001100000: M1r = 2'b01;
			14'b01001001100000: M1r = 2'b01;
			14'b10001001100000: M1r = 2'b10;
			14'b11001001100000: M1r = 2'b10;
			14'b00011001100000: M1r = 2'b01;
			14'b01011001100000: M1r = 2'b01;
			14'b10011001100000: M1r = 2'b01;
			14'b11011001100000: M1r = 2'b01;
			14'b00101001100000: M1r = 2'b00;
			14'b01101001100000: M1r = 2'b00;
			14'b10101001100000: M1r = 2'b01;
			14'b11101001100000: M1r = 2'b01;
			14'b00111001100000: M1r = 2'b00;
			14'b01111001100000: M1r = 2'b00;
			14'b10111001100000: M1r = 2'b00;
			14'b11111001100000: M1r = 2'b00;
			14'b00001101100000: M1r = 2'b10;
			14'b01001101100000: M1r = 2'b10;
			14'b10001101100000: M1r = 2'b10;
			14'b11001101100000: M1r = 2'b10;
			14'b00011101100000: M1r = 2'b01;
			14'b01011101100000: M1r = 2'b10;
			14'b10011101100000: M1r = 2'b10;
			14'b11011101100000: M1r = 2'b10;
			14'b00101101100000: M1r = 2'b01;
			14'b01101101100000: M1r = 2'b01;
			14'b10101101100000: M1r = 2'b01;
			14'b11101101100000: M1r = 2'b01;
			14'b00111101100000: M1r = 2'b01;
			14'b01111101100000: M1r = 2'b01;
			14'b10111101100000: M1r = 2'b01;
			14'b11111101100000: M1r = 2'b01;
			14'b00000010100000: M1r = 2'b00;
			14'b01000010100000: M1r = 2'b00;
			14'b10000010100000: M1r = 2'b00;
			14'b11000010100000: M1r = 2'b00;
			14'b00010010100000: M1r = 2'b00;
			14'b01010010100000: M1r = 2'b00;
			14'b10010010100000: M1r = 2'b00;
			14'b11010010100000: M1r = 2'b00;
			14'b00100010100000: M1r = 2'b00;
			14'b01100010100000: M1r = 2'b00;
			14'b10100010100000: M1r = 2'b00;
			14'b11100010100000: M1r = 2'b00;
			14'b00110010100000: M1r = 2'b00;
			14'b01110010100000: M1r = 2'b00;
			14'b10110010100000: M1r = 2'b00;
			14'b11110010100000: M1r = 2'b00;
			14'b00000110100000: M1r = 2'b00;
			14'b01000110100000: M1r = 2'b00;
			14'b10000110100000: M1r = 2'b01;
			14'b11000110100000: M1r = 2'b01;
			14'b00010110100000: M1r = 2'b00;
			14'b01010110100000: M1r = 2'b00;
			14'b10010110100000: M1r = 2'b00;
			14'b11010110100000: M1r = 2'b00;
			14'b00100110100000: M1r = 2'b00;
			14'b01100110100000: M1r = 2'b00;
			14'b10100110100000: M1r = 2'b00;
			14'b11100110100000: M1r = 2'b00;
			14'b00110110100000: M1r = 2'b00;
			14'b01110110100000: M1r = 2'b00;
			14'b10110110100000: M1r = 2'b00;
			14'b11110110100000: M1r = 2'b00;
			14'b00001010100000: M1r = 2'b01;
			14'b01001010100000: M1r = 2'b01;
			14'b10001010100000: M1r = 2'b01;
			14'b11001010100000: M1r = 2'b01;
			14'b00011010100000: M1r = 2'b00;
			14'b01011010100000: M1r = 2'b01;
			14'b10011010100000: M1r = 2'b01;
			14'b11011010100000: M1r = 2'b01;
			14'b00101010100000: M1r = 2'b00;
			14'b01101010100000: M1r = 2'b00;
			14'b10101010100000: M1r = 2'b00;
			14'b11101010100000: M1r = 2'b00;
			14'b00111010100000: M1r = 2'b00;
			14'b01111010100000: M1r = 2'b00;
			14'b10111010100000: M1r = 2'b00;
			14'b11111010100000: M1r = 2'b00;
			14'b00001110100000: M1r = 2'b10;
			14'b01001110100000: M1r = 2'b10;
			14'b10001110100000: M1r = 2'b10;
			14'b11001110100000: M1r = 2'b10;
			14'b00011110100000: M1r = 2'b01;
			14'b01011110100000: M1r = 2'b01;
			14'b10011110100000: M1r = 2'b10;
			14'b11011110100000: M1r = 2'b10;
			14'b00101110100000: M1r = 2'b01;
			14'b01101110100000: M1r = 2'b01;
			14'b10101110100000: M1r = 2'b01;
			14'b11101110100000: M1r = 2'b01;
			14'b00111110100000: M1r = 2'b00;
			14'b01111110100000: M1r = 2'b00;
			14'b10111110100000: M1r = 2'b01;
			14'b11111110100000: M1r = 2'b01;
			14'b00000011100000: M1r = 2'b00;
			14'b01000011100000: M1r = 2'b00;
			14'b10000011100000: M1r = 2'b00;
			14'b11000011100000: M1r = 2'b00;
			14'b00010011100000: M1r = 2'b00;
			14'b01010011100000: M1r = 2'b00;
			14'b10010011100000: M1r = 2'b00;
			14'b11010011100000: M1r = 2'b00;
			14'b00100011100000: M1r = 2'b00;
			14'b01100011100000: M1r = 2'b00;
			14'b10100011100000: M1r = 2'b00;
			14'b11100011100000: M1r = 2'b00;
			14'b00110011100000: M1r = 2'b00;
			14'b01110011100000: M1r = 2'b00;
			14'b10110011100000: M1r = 2'b00;
			14'b11110011100000: M1r = 2'b00;
			14'b00000111100000: M1r = 2'b00;
			14'b01000111100000: M1r = 2'b00;
			14'b10000111100000: M1r = 2'b00;
			14'b11000111100000: M1r = 2'b00;
			14'b00010111100000: M1r = 2'b00;
			14'b01010111100000: M1r = 2'b00;
			14'b10010111100000: M1r = 2'b00;
			14'b11010111100000: M1r = 2'b00;
			14'b00100111100000: M1r = 2'b00;
			14'b01100111100000: M1r = 2'b00;
			14'b10100111100000: M1r = 2'b00;
			14'b11100111100000: M1r = 2'b00;
			14'b00110111100000: M1r = 2'b00;
			14'b01110111100000: M1r = 2'b00;
			14'b10110111100000: M1r = 2'b00;
			14'b11110111100000: M1r = 2'b00;
			14'b00001011100000: M1r = 2'b01;
			14'b01001011100000: M1r = 2'b01;
			14'b10001011100000: M1r = 2'b01;
			14'b11001011100000: M1r = 2'b01;
			14'b00011011100000: M1r = 2'b00;
			14'b01011011100000: M1r = 2'b00;
			14'b10011011100000: M1r = 2'b01;
			14'b11011011100000: M1r = 2'b01;
			14'b00101011100000: M1r = 2'b00;
			14'b01101011100000: M1r = 2'b00;
			14'b10101011100000: M1r = 2'b00;
			14'b11101011100000: M1r = 2'b00;
			14'b00111011100000: M1r = 2'b00;
			14'b01111011100000: M1r = 2'b00;
			14'b10111011100000: M1r = 2'b00;
			14'b11111011100000: M1r = 2'b00;
			14'b00001111100000: M1r = 2'b01;
			14'b01001111100000: M1r = 2'b10;
			14'b10001111100000: M1r = 2'b10;
			14'b11001111100000: M1r = 2'b10;
			14'b00011111100000: M1r = 2'b01;
			14'b01011111100000: M1r = 2'b01;
			14'b10011111100000: M1r = 2'b01;
			14'b11011111100000: M1r = 2'b01;
			14'b00101111100000: M1r = 2'b00;
			14'b01101111100000: M1r = 2'b01;
			14'b10101111100000: M1r = 2'b01;
			14'b11101111100000: M1r = 2'b01;
			14'b00111111100000: M1r = 2'b00;
			14'b01111111100000: M1r = 2'b00;
			14'b10111111100000: M1r = 2'b00;
			14'b11111111100000: M1r = 2'b00;
			14'b00000000110000: M1r = 2'b00;
			14'b01000000110000: M1r = 2'b01;
			14'b10000000110000: M1r = 2'b01;
			14'b11000000110000: M1r = 2'b01;
			14'b00010000110000: M1r = 2'b00;
			14'b01010000110000: M1r = 2'b00;
			14'b10010000110000: M1r = 2'b00;
			14'b11010000110000: M1r = 2'b00;
			14'b00100000110000: M1r = 2'b00;
			14'b01100000110000: M1r = 2'b00;
			14'b10100000110000: M1r = 2'b00;
			14'b11100000110000: M1r = 2'b00;
			14'b00110000110000: M1r = 2'b00;
			14'b01110000110000: M1r = 2'b00;
			14'b10110000110000: M1r = 2'b00;
			14'b11110000110000: M1r = 2'b00;
			14'b00000100110000: M1r = 2'b01;
			14'b01000100110000: M1r = 2'b01;
			14'b10000100110000: M1r = 2'b01;
			14'b11000100110000: M1r = 2'b10;
			14'b00010100110000: M1r = 2'b01;
			14'b01010100110000: M1r = 2'b01;
			14'b10010100110000: M1r = 2'b01;
			14'b11010100110000: M1r = 2'b01;
			14'b00100100110000: M1r = 2'b00;
			14'b01100100110000: M1r = 2'b00;
			14'b10100100110000: M1r = 2'b01;
			14'b11100100110000: M1r = 2'b01;
			14'b00110100110000: M1r = 2'b00;
			14'b01110100110000: M1r = 2'b00;
			14'b10110100110000: M1r = 2'b00;
			14'b11110100110000: M1r = 2'b00;
			14'b00001000110000: M1r = 2'b10;
			14'b01001000110000: M1r = 2'b10;
			14'b10001000110000: M1r = 2'b10;
			14'b11001000110000: M1r = 2'b10;
			14'b00011000110000: M1r = 2'b01;
			14'b01011000110000: M1r = 2'b10;
			14'b10011000110000: M1r = 2'b10;
			14'b11011000110000: M1r = 2'b10;
			14'b00101000110000: M1r = 2'b01;
			14'b01101000110000: M1r = 2'b01;
			14'b10101000110000: M1r = 2'b01;
			14'b11101000110000: M1r = 2'b01;
			14'b00111000110000: M1r = 2'b01;
			14'b01111000110000: M1r = 2'b01;
			14'b10111000110000: M1r = 2'b01;
			14'b11111000110000: M1r = 2'b01;
			14'b00001100110000: M1r = 2'b11;
			14'b01001100110000: M1r = 2'b11;
			14'b10001100110000: M1r = 2'b11;
			14'b11001100110000: M1r = 2'b11;
			14'b00011100110000: M1r = 2'b10;
			14'b01011100110000: M1r = 2'b10;
			14'b10011100110000: M1r = 2'b11;
			14'b11011100110000: M1r = 2'b11;
			14'b00101100110000: M1r = 2'b10;
			14'b01101100110000: M1r = 2'b10;
			14'b10101100110000: M1r = 2'b10;
			14'b11101100110000: M1r = 2'b10;
			14'b00111100110000: M1r = 2'b01;
			14'b01111100110000: M1r = 2'b01;
			14'b10111100110000: M1r = 2'b10;
			14'b11111100110000: M1r = 2'b10;
			14'b00000001110000: M1r = 2'b00;
			14'b01000001110000: M1r = 2'b00;
			14'b10000001110000: M1r = 2'b00;
			14'b11000001110000: M1r = 2'b01;
			14'b00010001110000: M1r = 2'b00;
			14'b01010001110000: M1r = 2'b00;
			14'b10010001110000: M1r = 2'b00;
			14'b11010001110000: M1r = 2'b00;
			14'b00100001110000: M1r = 2'b00;
			14'b01100001110000: M1r = 2'b00;
			14'b10100001110000: M1r = 2'b00;
			14'b11100001110000: M1r = 2'b00;
			14'b00110001110000: M1r = 2'b00;
			14'b01110001110000: M1r = 2'b00;
			14'b10110001110000: M1r = 2'b00;
			14'b11110001110000: M1r = 2'b00;
			14'b00000101110000: M1r = 2'b01;
			14'b01000101110000: M1r = 2'b01;
			14'b10000101110000: M1r = 2'b01;
			14'b11000101110000: M1r = 2'b01;
			14'b00010101110000: M1r = 2'b00;
			14'b01010101110000: M1r = 2'b01;
			14'b10010101110000: M1r = 2'b01;
			14'b11010101110000: M1r = 2'b01;
			14'b00100101110000: M1r = 2'b00;
			14'b01100101110000: M1r = 2'b00;
			14'b10100101110000: M1r = 2'b00;
			14'b11100101110000: M1r = 2'b00;
			14'b00110101110000: M1r = 2'b00;
			14'b01110101110000: M1r = 2'b00;
			14'b10110101110000: M1r = 2'b00;
			14'b11110101110000: M1r = 2'b00;
			14'b00001001110000: M1r = 2'b10;
			14'b01001001110000: M1r = 2'b10;
			14'b10001001110000: M1r = 2'b10;
			14'b11001001110000: M1r = 2'b10;
			14'b00011001110000: M1r = 2'b01;
			14'b01011001110000: M1r = 2'b01;
			14'b10011001110000: M1r = 2'b01;
			14'b11011001110000: M1r = 2'b10;
			14'b00101001110000: M1r = 2'b01;
			14'b01101001110000: M1r = 2'b01;
			14'b10101001110000: M1r = 2'b01;
			14'b11101001110000: M1r = 2'b01;
			14'b00111001110000: M1r = 2'b00;
			14'b01111001110000: M1r = 2'b00;
			14'b10111001110000: M1r = 2'b01;
			14'b11111001110000: M1r = 2'b01;
			14'b00001101110000: M1r = 2'b10;
			14'b01001101110000: M1r = 2'b11;
			14'b10001101110000: M1r = 2'b11;
			14'b11001101110000: M1r = 2'b11;
			14'b00011101110000: M1r = 2'b10;
			14'b01011101110000: M1r = 2'b10;
			14'b10011101110000: M1r = 2'b10;
			14'b11011101110000: M1r = 2'b10;
			14'b00101101110000: M1r = 2'b01;
			14'b01101101110000: M1r = 2'b10;
			14'b10101101110000: M1r = 2'b10;
			14'b11101101110000: M1r = 2'b10;
			14'b00111101110000: M1r = 2'b01;
			14'b01111101110000: M1r = 2'b01;
			14'b10111101110000: M1r = 2'b01;
			14'b11111101110000: M1r = 2'b01;
			14'b00000010110000: M1r = 2'b00;
			14'b01000010110000: M1r = 2'b00;
			14'b10000010110000: M1r = 2'b00;
			14'b11000010110000: M1r = 2'b00;
			14'b00010010110000: M1r = 2'b00;
			14'b01010010110000: M1r = 2'b00;
			14'b10010010110000: M1r = 2'b00;
			14'b11010010110000: M1r = 2'b00;
			14'b00100010110000: M1r = 2'b00;
			14'b01100010110000: M1r = 2'b00;
			14'b10100010110000: M1r = 2'b00;
			14'b11100010110000: M1r = 2'b00;
			14'b00110010110000: M1r = 2'b00;
			14'b01110010110000: M1r = 2'b00;
			14'b10110010110000: M1r = 2'b00;
			14'b11110010110000: M1r = 2'b00;
			14'b00000110110000: M1r = 2'b01;
			14'b01000110110000: M1r = 2'b01;
			14'b10000110110000: M1r = 2'b01;
			14'b11000110110000: M1r = 2'b01;
			14'b00010110110000: M1r = 2'b00;
			14'b01010110110000: M1r = 2'b00;
			14'b10010110110000: M1r = 2'b00;
			14'b11010110110000: M1r = 2'b01;
			14'b00100110110000: M1r = 2'b00;
			14'b01100110110000: M1r = 2'b00;
			14'b10100110110000: M1r = 2'b00;
			14'b11100110110000: M1r = 2'b00;
			14'b00110110110000: M1r = 2'b00;
			14'b01110110110000: M1r = 2'b00;
			14'b10110110110000: M1r = 2'b00;
			14'b11110110110000: M1r = 2'b00;
			14'b00001010110000: M1r = 2'b01;
			14'b01001010110000: M1r = 2'b10;
			14'b10001010110000: M1r = 2'b10;
			14'b11001010110000: M1r = 2'b10;
			14'b00011010110000: M1r = 2'b01;
			14'b01011010110000: M1r = 2'b01;
			14'b10011010110000: M1r = 2'b01;
			14'b11011010110000: M1r = 2'b01;
			14'b00101010110000: M1r = 2'b00;
			14'b01101010110000: M1r = 2'b01;
			14'b10101010110000: M1r = 2'b01;
			14'b11101010110000: M1r = 2'b01;
			14'b00111010110000: M1r = 2'b00;
			14'b01111010110000: M1r = 2'b00;
			14'b10111010110000: M1r = 2'b00;
			14'b11111010110000: M1r = 2'b00;
			14'b00001110110000: M1r = 2'b10;
			14'b01001110110000: M1r = 2'b10;
			14'b10001110110000: M1r = 2'b10;
			14'b11001110110000: M1r = 2'b11;
			14'b00011110110000: M1r = 2'b10;
			14'b01011110110000: M1r = 2'b10;
			14'b10011110110000: M1r = 2'b10;
			14'b11011110110000: M1r = 2'b10;
			14'b00101110110000: M1r = 2'b01;
			14'b01101110110000: M1r = 2'b01;
			14'b10101110110000: M1r = 2'b01;
			14'b11101110110000: M1r = 2'b10;
			14'b00111110110000: M1r = 2'b01;
			14'b01111110110000: M1r = 2'b01;
			14'b10111110110000: M1r = 2'b01;
			14'b11111110110000: M1r = 2'b01;
			14'b00000011110000: M1r = 2'b00;
			14'b01000011110000: M1r = 2'b00;
			14'b10000011110000: M1r = 2'b00;
			14'b11000011110000: M1r = 2'b00;
			14'b00010011110000: M1r = 2'b00;
			14'b01010011110000: M1r = 2'b00;
			14'b10010011110000: M1r = 2'b00;
			14'b11010011110000: M1r = 2'b00;
			14'b00100011110000: M1r = 2'b00;
			14'b01100011110000: M1r = 2'b00;
			14'b10100011110000: M1r = 2'b00;
			14'b11100011110000: M1r = 2'b00;
			14'b00110011110000: M1r = 2'b00;
			14'b01110011110000: M1r = 2'b00;
			14'b10110011110000: M1r = 2'b00;
			14'b11110011110000: M1r = 2'b00;
			14'b00000111110000: M1r = 2'b00;
			14'b01000111110000: M1r = 2'b01;
			14'b10000111110000: M1r = 2'b01;
			14'b11000111110000: M1r = 2'b01;
			14'b00010111110000: M1r = 2'b00;
			14'b01010111110000: M1r = 2'b00;
			14'b10010111110000: M1r = 2'b00;
			14'b11010111110000: M1r = 2'b00;
			14'b00100111110000: M1r = 2'b00;
			14'b01100111110000: M1r = 2'b00;
			14'b10100111110000: M1r = 2'b00;
			14'b11100111110000: M1r = 2'b00;
			14'b00110111110000: M1r = 2'b00;
			14'b01110111110000: M1r = 2'b00;
			14'b10110111110000: M1r = 2'b00;
			14'b11110111110000: M1r = 2'b00;
			14'b00001011110000: M1r = 2'b01;
			14'b01001011110000: M1r = 2'b01;
			14'b10001011110000: M1r = 2'b01;
			14'b11001011110000: M1r = 2'b10;
			14'b00011011110000: M1r = 2'b01;
			14'b01011011110000: M1r = 2'b01;
			14'b10011011110000: M1r = 2'b01;
			14'b11011011110000: M1r = 2'b01;
			14'b00101011110000: M1r = 2'b00;
			14'b01101011110000: M1r = 2'b00;
			14'b10101011110000: M1r = 2'b00;
			14'b11101011110000: M1r = 2'b01;
			14'b00111011110000: M1r = 2'b00;
			14'b01111011110000: M1r = 2'b00;
			14'b10111011110000: M1r = 2'b00;
			14'b11111011110000: M1r = 2'b00;
			14'b00001111110000: M1r = 2'b10;
			14'b01001111110000: M1r = 2'b10;
			14'b10001111110000: M1r = 2'b10;
			14'b11001111110000: M1r = 2'b10;
			14'b00011111110000: M1r = 2'b01;
			14'b01011111110000: M1r = 2'b10;
			14'b10011111110000: M1r = 2'b10;
			14'b11011111110000: M1r = 2'b10;
			14'b00101111110000: M1r = 2'b01;
			14'b01101111110000: M1r = 2'b01;
			14'b10101111110000: M1r = 2'b01;
			14'b11101111110000: M1r = 2'b01;
			14'b00111111110000: M1r = 2'b00;
			14'b01111111110000: M1r = 2'b01;
			14'b10111111110000: M1r = 2'b01;
			14'b11111111110000: M1r = 2'b01;
			14'b00000000000100: M1r = 2'b00;
			14'b01000000000100: M1r = 2'b00;
			14'b10000000000100: M1r = 2'b00;
			14'b11000000000100: M1r = 2'b00;
			14'b00010000000100: M1r = 2'b00;
			14'b01010000000100: M1r = 2'b00;
			14'b10010000000100: M1r = 2'b00;
			14'b11010000000100: M1r = 2'b00;
			14'b00100000000100: M1r = 2'b00;
			14'b01100000000100: M1r = 2'b00;
			14'b10100000000100: M1r = 2'b00;
			14'b11100000000100: M1r = 2'b00;
			14'b00110000000100: M1r = 2'b00;
			14'b01110000000100: M1r = 2'b00;
			14'b10110000000100: M1r = 2'b00;
			14'b11110000000100: M1r = 2'b00;
			14'b00000100000100: M1r = 2'b00;
			14'b01000100000100: M1r = 2'b00;
			14'b10000100000100: M1r = 2'b00;
			14'b11000100000100: M1r = 2'b00;
			14'b00010100000100: M1r = 2'b00;
			14'b01010100000100: M1r = 2'b00;
			14'b10010100000100: M1r = 2'b00;
			14'b11010100000100: M1r = 2'b00;
			14'b00100100000100: M1r = 2'b00;
			14'b01100100000100: M1r = 2'b00;
			14'b10100100000100: M1r = 2'b00;
			14'b11100100000100: M1r = 2'b00;
			14'b00110100000100: M1r = 2'b00;
			14'b01110100000100: M1r = 2'b00;
			14'b10110100000100: M1r = 2'b00;
			14'b11110100000100: M1r = 2'b00;
			14'b00001000000100: M1r = 2'b00;
			14'b01001000000100: M1r = 2'b00;
			14'b10001000000100: M1r = 2'b00;
			14'b11001000000100: M1r = 2'b00;
			14'b00011000000100: M1r = 2'b00;
			14'b01011000000100: M1r = 2'b00;
			14'b10011000000100: M1r = 2'b00;
			14'b11011000000100: M1r = 2'b00;
			14'b00101000000100: M1r = 2'b00;
			14'b01101000000100: M1r = 2'b00;
			14'b10101000000100: M1r = 2'b00;
			14'b11101000000100: M1r = 2'b00;
			14'b00111000000100: M1r = 2'b00;
			14'b01111000000100: M1r = 2'b00;
			14'b10111000000100: M1r = 2'b00;
			14'b11111000000100: M1r = 2'b00;
			14'b00001100000100: M1r = 2'b01;
			14'b01001100000100: M1r = 2'b01;
			14'b10001100000100: M1r = 2'b01;
			14'b11001100000100: M1r = 2'b01;
			14'b00011100000100: M1r = 2'b00;
			14'b01011100000100: M1r = 2'b00;
			14'b10011100000100: M1r = 2'b00;
			14'b11011100000100: M1r = 2'b01;
			14'b00101100000100: M1r = 2'b00;
			14'b01101100000100: M1r = 2'b00;
			14'b10101100000100: M1r = 2'b00;
			14'b11101100000100: M1r = 2'b00;
			14'b00111100000100: M1r = 2'b00;
			14'b01111100000100: M1r = 2'b00;
			14'b10111100000100: M1r = 2'b00;
			14'b11111100000100: M1r = 2'b00;
			14'b00000001000100: M1r = 2'b00;
			14'b01000001000100: M1r = 2'b00;
			14'b10000001000100: M1r = 2'b00;
			14'b11000001000100: M1r = 2'b00;
			14'b00010001000100: M1r = 2'b00;
			14'b01010001000100: M1r = 2'b00;
			14'b10010001000100: M1r = 2'b00;
			14'b11010001000100: M1r = 2'b00;
			14'b00100001000100: M1r = 2'b00;
			14'b01100001000100: M1r = 2'b00;
			14'b10100001000100: M1r = 2'b00;
			14'b11100001000100: M1r = 2'b00;
			14'b00110001000100: M1r = 2'b00;
			14'b01110001000100: M1r = 2'b00;
			14'b10110001000100: M1r = 2'b00;
			14'b11110001000100: M1r = 2'b00;
			14'b00000101000100: M1r = 2'b00;
			14'b01000101000100: M1r = 2'b00;
			14'b10000101000100: M1r = 2'b00;
			14'b11000101000100: M1r = 2'b00;
			14'b00010101000100: M1r = 2'b00;
			14'b01010101000100: M1r = 2'b00;
			14'b10010101000100: M1r = 2'b00;
			14'b11010101000100: M1r = 2'b00;
			14'b00100101000100: M1r = 2'b00;
			14'b01100101000100: M1r = 2'b00;
			14'b10100101000100: M1r = 2'b00;
			14'b11100101000100: M1r = 2'b00;
			14'b00110101000100: M1r = 2'b00;
			14'b01110101000100: M1r = 2'b00;
			14'b10110101000100: M1r = 2'b00;
			14'b11110101000100: M1r = 2'b00;
			14'b00001001000100: M1r = 2'b00;
			14'b01001001000100: M1r = 2'b00;
			14'b10001001000100: M1r = 2'b00;
			14'b11001001000100: M1r = 2'b00;
			14'b00011001000100: M1r = 2'b00;
			14'b01011001000100: M1r = 2'b00;
			14'b10011001000100: M1r = 2'b00;
			14'b11011001000100: M1r = 2'b00;
			14'b00101001000100: M1r = 2'b00;
			14'b01101001000100: M1r = 2'b00;
			14'b10101001000100: M1r = 2'b00;
			14'b11101001000100: M1r = 2'b00;
			14'b00111001000100: M1r = 2'b00;
			14'b01111001000100: M1r = 2'b00;
			14'b10111001000100: M1r = 2'b00;
			14'b11111001000100: M1r = 2'b00;
			14'b00001101000100: M1r = 2'b00;
			14'b01001101000100: M1r = 2'b00;
			14'b10001101000100: M1r = 2'b01;
			14'b11001101000100: M1r = 2'b01;
			14'b00011101000100: M1r = 2'b00;
			14'b01011101000100: M1r = 2'b00;
			14'b10011101000100: M1r = 2'b00;
			14'b11011101000100: M1r = 2'b00;
			14'b00101101000100: M1r = 2'b00;
			14'b01101101000100: M1r = 2'b00;
			14'b10101101000100: M1r = 2'b00;
			14'b11101101000100: M1r = 2'b00;
			14'b00111101000100: M1r = 2'b00;
			14'b01111101000100: M1r = 2'b00;
			14'b10111101000100: M1r = 2'b00;
			14'b11111101000100: M1r = 2'b00;
			14'b00000010000100: M1r = 2'b00;
			14'b01000010000100: M1r = 2'b00;
			14'b10000010000100: M1r = 2'b00;
			14'b11000010000100: M1r = 2'b00;
			14'b00010010000100: M1r = 2'b00;
			14'b01010010000100: M1r = 2'b00;
			14'b10010010000100: M1r = 2'b00;
			14'b11010010000100: M1r = 2'b00;
			14'b00100010000100: M1r = 2'b00;
			14'b01100010000100: M1r = 2'b00;
			14'b10100010000100: M1r = 2'b00;
			14'b11100010000100: M1r = 2'b00;
			14'b00110010000100: M1r = 2'b00;
			14'b01110010000100: M1r = 2'b00;
			14'b10110010000100: M1r = 2'b00;
			14'b11110010000100: M1r = 2'b00;
			14'b00000110000100: M1r = 2'b00;
			14'b01000110000100: M1r = 2'b00;
			14'b10000110000100: M1r = 2'b00;
			14'b11000110000100: M1r = 2'b00;
			14'b00010110000100: M1r = 2'b00;
			14'b01010110000100: M1r = 2'b00;
			14'b10010110000100: M1r = 2'b00;
			14'b11010110000100: M1r = 2'b00;
			14'b00100110000100: M1r = 2'b00;
			14'b01100110000100: M1r = 2'b00;
			14'b10100110000100: M1r = 2'b00;
			14'b11100110000100: M1r = 2'b00;
			14'b00110110000100: M1r = 2'b00;
			14'b01110110000100: M1r = 2'b00;
			14'b10110110000100: M1r = 2'b00;
			14'b11110110000100: M1r = 2'b00;
			14'b00001010000100: M1r = 2'b00;
			14'b01001010000100: M1r = 2'b00;
			14'b10001010000100: M1r = 2'b00;
			14'b11001010000100: M1r = 2'b00;
			14'b00011010000100: M1r = 2'b00;
			14'b01011010000100: M1r = 2'b00;
			14'b10011010000100: M1r = 2'b00;
			14'b11011010000100: M1r = 2'b00;
			14'b00101010000100: M1r = 2'b00;
			14'b01101010000100: M1r = 2'b00;
			14'b10101010000100: M1r = 2'b00;
			14'b11101010000100: M1r = 2'b00;
			14'b00111010000100: M1r = 2'b00;
			14'b01111010000100: M1r = 2'b00;
			14'b10111010000100: M1r = 2'b00;
			14'b11111010000100: M1r = 2'b00;
			14'b00001110000100: M1r = 2'b00;
			14'b01001110000100: M1r = 2'b00;
			14'b10001110000100: M1r = 2'b00;
			14'b11001110000100: M1r = 2'b01;
			14'b00011110000100: M1r = 2'b00;
			14'b01011110000100: M1r = 2'b00;
			14'b10011110000100: M1r = 2'b00;
			14'b11011110000100: M1r = 2'b00;
			14'b00101110000100: M1r = 2'b00;
			14'b01101110000100: M1r = 2'b00;
			14'b10101110000100: M1r = 2'b00;
			14'b11101110000100: M1r = 2'b00;
			14'b00111110000100: M1r = 2'b00;
			14'b01111110000100: M1r = 2'b00;
			14'b10111110000100: M1r = 2'b00;
			14'b11111110000100: M1r = 2'b00;
			14'b00000011000100: M1r = 2'b00;
			14'b01000011000100: M1r = 2'b00;
			14'b10000011000100: M1r = 2'b00;
			14'b11000011000100: M1r = 2'b00;
			14'b00010011000100: M1r = 2'b00;
			14'b01010011000100: M1r = 2'b00;
			14'b10010011000100: M1r = 2'b00;
			14'b11010011000100: M1r = 2'b00;
			14'b00100011000100: M1r = 2'b00;
			14'b01100011000100: M1r = 2'b00;
			14'b10100011000100: M1r = 2'b00;
			14'b11100011000100: M1r = 2'b00;
			14'b00110011000100: M1r = 2'b00;
			14'b01110011000100: M1r = 2'b00;
			14'b10110011000100: M1r = 2'b00;
			14'b11110011000100: M1r = 2'b00;
			14'b00000111000100: M1r = 2'b00;
			14'b01000111000100: M1r = 2'b00;
			14'b10000111000100: M1r = 2'b00;
			14'b11000111000100: M1r = 2'b00;
			14'b00010111000100: M1r = 2'b00;
			14'b01010111000100: M1r = 2'b00;
			14'b10010111000100: M1r = 2'b00;
			14'b11010111000100: M1r = 2'b00;
			14'b00100111000100: M1r = 2'b00;
			14'b01100111000100: M1r = 2'b00;
			14'b10100111000100: M1r = 2'b00;
			14'b11100111000100: M1r = 2'b00;
			14'b00110111000100: M1r = 2'b00;
			14'b01110111000100: M1r = 2'b00;
			14'b10110111000100: M1r = 2'b00;
			14'b11110111000100: M1r = 2'b00;
			14'b00001011000100: M1r = 2'b00;
			14'b01001011000100: M1r = 2'b00;
			14'b10001011000100: M1r = 2'b00;
			14'b11001011000100: M1r = 2'b00;
			14'b00011011000100: M1r = 2'b00;
			14'b01011011000100: M1r = 2'b00;
			14'b10011011000100: M1r = 2'b00;
			14'b11011011000100: M1r = 2'b00;
			14'b00101011000100: M1r = 2'b00;
			14'b01101011000100: M1r = 2'b00;
			14'b10101011000100: M1r = 2'b00;
			14'b11101011000100: M1r = 2'b00;
			14'b00111011000100: M1r = 2'b00;
			14'b01111011000100: M1r = 2'b00;
			14'b10111011000100: M1r = 2'b00;
			14'b11111011000100: M1r = 2'b00;
			14'b00001111000100: M1r = 2'b00;
			14'b01001111000100: M1r = 2'b00;
			14'b10001111000100: M1r = 2'b00;
			14'b11001111000100: M1r = 2'b00;
			14'b00011111000100: M1r = 2'b00;
			14'b01011111000100: M1r = 2'b00;
			14'b10011111000100: M1r = 2'b00;
			14'b11011111000100: M1r = 2'b00;
			14'b00101111000100: M1r = 2'b00;
			14'b01101111000100: M1r = 2'b00;
			14'b10101111000100: M1r = 2'b00;
			14'b11101111000100: M1r = 2'b00;
			14'b00111111000100: M1r = 2'b00;
			14'b01111111000100: M1r = 2'b00;
			14'b10111111000100: M1r = 2'b00;
			14'b11111111000100: M1r = 2'b00;
			14'b00000000010100: M1r = 2'b00;
			14'b01000000010100: M1r = 2'b00;
			14'b10000000010100: M1r = 2'b00;
			14'b11000000010100: M1r = 2'b00;
			14'b00010000010100: M1r = 2'b00;
			14'b01010000010100: M1r = 2'b00;
			14'b10010000010100: M1r = 2'b00;
			14'b11010000010100: M1r = 2'b00;
			14'b00100000010100: M1r = 2'b00;
			14'b01100000010100: M1r = 2'b00;
			14'b10100000010100: M1r = 2'b00;
			14'b11100000010100: M1r = 2'b00;
			14'b00110000010100: M1r = 2'b00;
			14'b01110000010100: M1r = 2'b00;
			14'b10110000010100: M1r = 2'b00;
			14'b11110000010100: M1r = 2'b00;
			14'b00000100010100: M1r = 2'b00;
			14'b01000100010100: M1r = 2'b00;
			14'b10000100010100: M1r = 2'b00;
			14'b11000100010100: M1r = 2'b00;
			14'b00010100010100: M1r = 2'b00;
			14'b01010100010100: M1r = 2'b00;
			14'b10010100010100: M1r = 2'b00;
			14'b11010100010100: M1r = 2'b00;
			14'b00100100010100: M1r = 2'b00;
			14'b01100100010100: M1r = 2'b00;
			14'b10100100010100: M1r = 2'b00;
			14'b11100100010100: M1r = 2'b00;
			14'b00110100010100: M1r = 2'b00;
			14'b01110100010100: M1r = 2'b00;
			14'b10110100010100: M1r = 2'b00;
			14'b11110100010100: M1r = 2'b00;
			14'b00001000010100: M1r = 2'b00;
			14'b01001000010100: M1r = 2'b00;
			14'b10001000010100: M1r = 2'b01;
			14'b11001000010100: M1r = 2'b01;
			14'b00011000010100: M1r = 2'b00;
			14'b01011000010100: M1r = 2'b00;
			14'b10011000010100: M1r = 2'b00;
			14'b11011000010100: M1r = 2'b00;
			14'b00101000010100: M1r = 2'b00;
			14'b01101000010100: M1r = 2'b00;
			14'b10101000010100: M1r = 2'b00;
			14'b11101000010100: M1r = 2'b00;
			14'b00111000010100: M1r = 2'b00;
			14'b01111000010100: M1r = 2'b00;
			14'b10111000010100: M1r = 2'b00;
			14'b11111000010100: M1r = 2'b00;
			14'b00001100010100: M1r = 2'b01;
			14'b01001100010100: M1r = 2'b01;
			14'b10001100010100: M1r = 2'b01;
			14'b11001100010100: M1r = 2'b01;
			14'b00011100010100: M1r = 2'b01;
			14'b01011100010100: M1r = 2'b01;
			14'b10011100010100: M1r = 2'b01;
			14'b11011100010100: M1r = 2'b01;
			14'b00101100010100: M1r = 2'b00;
			14'b01101100010100: M1r = 2'b00;
			14'b10101100010100: M1r = 2'b00;
			14'b11101100010100: M1r = 2'b01;
			14'b00111100010100: M1r = 2'b00;
			14'b01111100010100: M1r = 2'b00;
			14'b10111100010100: M1r = 2'b00;
			14'b11111100010100: M1r = 2'b00;
			14'b00000001010100: M1r = 2'b00;
			14'b01000001010100: M1r = 2'b00;
			14'b10000001010100: M1r = 2'b00;
			14'b11000001010100: M1r = 2'b00;
			14'b00010001010100: M1r = 2'b00;
			14'b01010001010100: M1r = 2'b00;
			14'b10010001010100: M1r = 2'b00;
			14'b11010001010100: M1r = 2'b00;
			14'b00100001010100: M1r = 2'b00;
			14'b01100001010100: M1r = 2'b00;
			14'b10100001010100: M1r = 2'b00;
			14'b11100001010100: M1r = 2'b00;
			14'b00110001010100: M1r = 2'b00;
			14'b01110001010100: M1r = 2'b00;
			14'b10110001010100: M1r = 2'b00;
			14'b11110001010100: M1r = 2'b00;
			14'b00000101010100: M1r = 2'b00;
			14'b01000101010100: M1r = 2'b00;
			14'b10000101010100: M1r = 2'b00;
			14'b11000101010100: M1r = 2'b00;
			14'b00010101010100: M1r = 2'b00;
			14'b01010101010100: M1r = 2'b00;
			14'b10010101010100: M1r = 2'b00;
			14'b11010101010100: M1r = 2'b00;
			14'b00100101010100: M1r = 2'b00;
			14'b01100101010100: M1r = 2'b00;
			14'b10100101010100: M1r = 2'b00;
			14'b11100101010100: M1r = 2'b00;
			14'b00110101010100: M1r = 2'b00;
			14'b01110101010100: M1r = 2'b00;
			14'b10110101010100: M1r = 2'b00;
			14'b11110101010100: M1r = 2'b00;
			14'b00001001010100: M1r = 2'b00;
			14'b01001001010100: M1r = 2'b00;
			14'b10001001010100: M1r = 2'b00;
			14'b11001001010100: M1r = 2'b00;
			14'b00011001010100: M1r = 2'b00;
			14'b01011001010100: M1r = 2'b00;
			14'b10011001010100: M1r = 2'b00;
			14'b11011001010100: M1r = 2'b00;
			14'b00101001010100: M1r = 2'b00;
			14'b01101001010100: M1r = 2'b00;
			14'b10101001010100: M1r = 2'b00;
			14'b11101001010100: M1r = 2'b00;
			14'b00111001010100: M1r = 2'b00;
			14'b01111001010100: M1r = 2'b00;
			14'b10111001010100: M1r = 2'b00;
			14'b11111001010100: M1r = 2'b00;
			14'b00001101010100: M1r = 2'b01;
			14'b01001101010100: M1r = 2'b01;
			14'b10001101010100: M1r = 2'b01;
			14'b11001101010100: M1r = 2'b01;
			14'b00011101010100: M1r = 2'b00;
			14'b01011101010100: M1r = 2'b00;
			14'b10011101010100: M1r = 2'b01;
			14'b11011101010100: M1r = 2'b01;
			14'b00101101010100: M1r = 2'b00;
			14'b01101101010100: M1r = 2'b00;
			14'b10101101010100: M1r = 2'b00;
			14'b11101101010100: M1r = 2'b00;
			14'b00111101010100: M1r = 2'b00;
			14'b01111101010100: M1r = 2'b00;
			14'b10111101010100: M1r = 2'b00;
			14'b11111101010100: M1r = 2'b00;
			14'b00000010010100: M1r = 2'b00;
			14'b01000010010100: M1r = 2'b00;
			14'b10000010010100: M1r = 2'b00;
			14'b11000010010100: M1r = 2'b00;
			14'b00010010010100: M1r = 2'b00;
			14'b01010010010100: M1r = 2'b00;
			14'b10010010010100: M1r = 2'b00;
			14'b11010010010100: M1r = 2'b00;
			14'b00100010010100: M1r = 2'b00;
			14'b01100010010100: M1r = 2'b00;
			14'b10100010010100: M1r = 2'b00;
			14'b11100010010100: M1r = 2'b00;
			14'b00110010010100: M1r = 2'b00;
			14'b01110010010100: M1r = 2'b00;
			14'b10110010010100: M1r = 2'b00;
			14'b11110010010100: M1r = 2'b00;
			14'b00000110010100: M1r = 2'b00;
			14'b01000110010100: M1r = 2'b00;
			14'b10000110010100: M1r = 2'b00;
			14'b11000110010100: M1r = 2'b00;
			14'b00010110010100: M1r = 2'b00;
			14'b01010110010100: M1r = 2'b00;
			14'b10010110010100: M1r = 2'b00;
			14'b11010110010100: M1r = 2'b00;
			14'b00100110010100: M1r = 2'b00;
			14'b01100110010100: M1r = 2'b00;
			14'b10100110010100: M1r = 2'b00;
			14'b11100110010100: M1r = 2'b00;
			14'b00110110010100: M1r = 2'b00;
			14'b01110110010100: M1r = 2'b00;
			14'b10110110010100: M1r = 2'b00;
			14'b11110110010100: M1r = 2'b00;
			14'b00001010010100: M1r = 2'b00;
			14'b01001010010100: M1r = 2'b00;
			14'b10001010010100: M1r = 2'b00;
			14'b11001010010100: M1r = 2'b00;
			14'b00011010010100: M1r = 2'b00;
			14'b01011010010100: M1r = 2'b00;
			14'b10011010010100: M1r = 2'b00;
			14'b11011010010100: M1r = 2'b00;
			14'b00101010010100: M1r = 2'b00;
			14'b01101010010100: M1r = 2'b00;
			14'b10101010010100: M1r = 2'b00;
			14'b11101010010100: M1r = 2'b00;
			14'b00111010010100: M1r = 2'b00;
			14'b01111010010100: M1r = 2'b00;
			14'b10111010010100: M1r = 2'b00;
			14'b11111010010100: M1r = 2'b00;
			14'b00001110010100: M1r = 2'b00;
			14'b01001110010100: M1r = 2'b01;
			14'b10001110010100: M1r = 2'b01;
			14'b11001110010100: M1r = 2'b01;
			14'b00011110010100: M1r = 2'b00;
			14'b01011110010100: M1r = 2'b00;
			14'b10011110010100: M1r = 2'b00;
			14'b11011110010100: M1r = 2'b00;
			14'b00101110010100: M1r = 2'b00;
			14'b01101110010100: M1r = 2'b00;
			14'b10101110010100: M1r = 2'b00;
			14'b11101110010100: M1r = 2'b00;
			14'b00111110010100: M1r = 2'b00;
			14'b01111110010100: M1r = 2'b00;
			14'b10111110010100: M1r = 2'b00;
			14'b11111110010100: M1r = 2'b00;
			14'b00000011010100: M1r = 2'b00;
			14'b01000011010100: M1r = 2'b00;
			14'b10000011010100: M1r = 2'b00;
			14'b11000011010100: M1r = 2'b00;
			14'b00010011010100: M1r = 2'b00;
			14'b01010011010100: M1r = 2'b00;
			14'b10010011010100: M1r = 2'b00;
			14'b11010011010100: M1r = 2'b00;
			14'b00100011010100: M1r = 2'b00;
			14'b01100011010100: M1r = 2'b00;
			14'b10100011010100: M1r = 2'b00;
			14'b11100011010100: M1r = 2'b00;
			14'b00110011010100: M1r = 2'b00;
			14'b01110011010100: M1r = 2'b00;
			14'b10110011010100: M1r = 2'b00;
			14'b11110011010100: M1r = 2'b00;
			14'b00000111010100: M1r = 2'b00;
			14'b01000111010100: M1r = 2'b00;
			14'b10000111010100: M1r = 2'b00;
			14'b11000111010100: M1r = 2'b00;
			14'b00010111010100: M1r = 2'b00;
			14'b01010111010100: M1r = 2'b00;
			14'b10010111010100: M1r = 2'b00;
			14'b11010111010100: M1r = 2'b00;
			14'b00100111010100: M1r = 2'b00;
			14'b01100111010100: M1r = 2'b00;
			14'b10100111010100: M1r = 2'b00;
			14'b11100111010100: M1r = 2'b00;
			14'b00110111010100: M1r = 2'b00;
			14'b01110111010100: M1r = 2'b00;
			14'b10110111010100: M1r = 2'b00;
			14'b11110111010100: M1r = 2'b00;
			14'b00001011010100: M1r = 2'b00;
			14'b01001011010100: M1r = 2'b00;
			14'b10001011010100: M1r = 2'b00;
			14'b11001011010100: M1r = 2'b00;
			14'b00011011010100: M1r = 2'b00;
			14'b01011011010100: M1r = 2'b00;
			14'b10011011010100: M1r = 2'b00;
			14'b11011011010100: M1r = 2'b00;
			14'b00101011010100: M1r = 2'b00;
			14'b01101011010100: M1r = 2'b00;
			14'b10101011010100: M1r = 2'b00;
			14'b11101011010100: M1r = 2'b00;
			14'b00111011010100: M1r = 2'b00;
			14'b01111011010100: M1r = 2'b00;
			14'b10111011010100: M1r = 2'b00;
			14'b11111011010100: M1r = 2'b00;
			14'b00001111010100: M1r = 2'b00;
			14'b01001111010100: M1r = 2'b00;
			14'b10001111010100: M1r = 2'b01;
			14'b11001111010100: M1r = 2'b01;
			14'b00011111010100: M1r = 2'b00;
			14'b01011111010100: M1r = 2'b00;
			14'b10011111010100: M1r = 2'b00;
			14'b11011111010100: M1r = 2'b00;
			14'b00101111010100: M1r = 2'b00;
			14'b01101111010100: M1r = 2'b00;
			14'b10101111010100: M1r = 2'b00;
			14'b11101111010100: M1r = 2'b00;
			14'b00111111010100: M1r = 2'b00;
			14'b01111111010100: M1r = 2'b00;
			14'b10111111010100: M1r = 2'b00;
			14'b11111111010100: M1r = 2'b00;
			14'b00000000100100: M1r = 2'b00;
			14'b01000000100100: M1r = 2'b00;
			14'b10000000100100: M1r = 2'b00;
			14'b11000000100100: M1r = 2'b00;
			14'b00010000100100: M1r = 2'b00;
			14'b01010000100100: M1r = 2'b00;
			14'b10010000100100: M1r = 2'b00;
			14'b11010000100100: M1r = 2'b00;
			14'b00100000100100: M1r = 2'b00;
			14'b01100000100100: M1r = 2'b00;
			14'b10100000100100: M1r = 2'b00;
			14'b11100000100100: M1r = 2'b00;
			14'b00110000100100: M1r = 2'b00;
			14'b01110000100100: M1r = 2'b00;
			14'b10110000100100: M1r = 2'b00;
			14'b11110000100100: M1r = 2'b00;
			14'b00000100100100: M1r = 2'b00;
			14'b01000100100100: M1r = 2'b00;
			14'b10000100100100: M1r = 2'b00;
			14'b11000100100100: M1r = 2'b00;
			14'b00010100100100: M1r = 2'b00;
			14'b01010100100100: M1r = 2'b00;
			14'b10010100100100: M1r = 2'b00;
			14'b11010100100100: M1r = 2'b00;
			14'b00100100100100: M1r = 2'b00;
			14'b01100100100100: M1r = 2'b00;
			14'b10100100100100: M1r = 2'b00;
			14'b11100100100100: M1r = 2'b00;
			14'b00110100100100: M1r = 2'b00;
			14'b01110100100100: M1r = 2'b00;
			14'b10110100100100: M1r = 2'b00;
			14'b11110100100100: M1r = 2'b00;
			14'b00001000100100: M1r = 2'b01;
			14'b01001000100100: M1r = 2'b01;
			14'b10001000100100: M1r = 2'b01;
			14'b11001000100100: M1r = 2'b01;
			14'b00011000100100: M1r = 2'b00;
			14'b01011000100100: M1r = 2'b00;
			14'b10011000100100: M1r = 2'b01;
			14'b11011000100100: M1r = 2'b01;
			14'b00101000100100: M1r = 2'b00;
			14'b01101000100100: M1r = 2'b00;
			14'b10101000100100: M1r = 2'b00;
			14'b11101000100100: M1r = 2'b00;
			14'b00111000100100: M1r = 2'b00;
			14'b01111000100100: M1r = 2'b00;
			14'b10111000100100: M1r = 2'b00;
			14'b11111000100100: M1r = 2'b00;
			14'b00001100100100: M1r = 2'b01;
			14'b01001100100100: M1r = 2'b10;
			14'b10001100100100: M1r = 2'b10;
			14'b11001100100100: M1r = 2'b10;
			14'b00011100100100: M1r = 2'b01;
			14'b01011100100100: M1r = 2'b01;
			14'b10011100100100: M1r = 2'b01;
			14'b11011100100100: M1r = 2'b01;
			14'b00101100100100: M1r = 2'b01;
			14'b01101100100100: M1r = 2'b01;
			14'b10101100100100: M1r = 2'b01;
			14'b11101100100100: M1r = 2'b01;
			14'b00111100100100: M1r = 2'b00;
			14'b01111100100100: M1r = 2'b00;
			14'b10111100100100: M1r = 2'b00;
			14'b11111100100100: M1r = 2'b01;
			14'b00000001100100: M1r = 2'b00;
			14'b01000001100100: M1r = 2'b00;
			14'b10000001100100: M1r = 2'b00;
			14'b11000001100100: M1r = 2'b00;
			14'b00010001100100: M1r = 2'b00;
			14'b01010001100100: M1r = 2'b00;
			14'b10010001100100: M1r = 2'b00;
			14'b11010001100100: M1r = 2'b00;
			14'b00100001100100: M1r = 2'b00;
			14'b01100001100100: M1r = 2'b00;
			14'b10100001100100: M1r = 2'b00;
			14'b11100001100100: M1r = 2'b00;
			14'b00110001100100: M1r = 2'b00;
			14'b01110001100100: M1r = 2'b00;
			14'b10110001100100: M1r = 2'b00;
			14'b11110001100100: M1r = 2'b00;
			14'b00000101100100: M1r = 2'b00;
			14'b01000101100100: M1r = 2'b00;
			14'b10000101100100: M1r = 2'b00;
			14'b11000101100100: M1r = 2'b00;
			14'b00010101100100: M1r = 2'b00;
			14'b01010101100100: M1r = 2'b00;
			14'b10010101100100: M1r = 2'b00;
			14'b11010101100100: M1r = 2'b00;
			14'b00100101100100: M1r = 2'b00;
			14'b01100101100100: M1r = 2'b00;
			14'b10100101100100: M1r = 2'b00;
			14'b11100101100100: M1r = 2'b00;
			14'b00110101100100: M1r = 2'b00;
			14'b01110101100100: M1r = 2'b00;
			14'b10110101100100: M1r = 2'b00;
			14'b11110101100100: M1r = 2'b00;
			14'b00001001100100: M1r = 2'b00;
			14'b01001001100100: M1r = 2'b01;
			14'b10001001100100: M1r = 2'b01;
			14'b11001001100100: M1r = 2'b01;
			14'b00011001100100: M1r = 2'b00;
			14'b01011001100100: M1r = 2'b00;
			14'b10011001100100: M1r = 2'b00;
			14'b11011001100100: M1r = 2'b00;
			14'b00101001100100: M1r = 2'b00;
			14'b01101001100100: M1r = 2'b00;
			14'b10101001100100: M1r = 2'b00;
			14'b11101001100100: M1r = 2'b00;
			14'b00111001100100: M1r = 2'b00;
			14'b01111001100100: M1r = 2'b00;
			14'b10111001100100: M1r = 2'b00;
			14'b11111001100100: M1r = 2'b00;
			14'b00001101100100: M1r = 2'b01;
			14'b01001101100100: M1r = 2'b01;
			14'b10001101100100: M1r = 2'b10;
			14'b11001101100100: M1r = 2'b10;
			14'b00011101100100: M1r = 2'b01;
			14'b01011101100100: M1r = 2'b01;
			14'b10011101100100: M1r = 2'b01;
			14'b11011101100100: M1r = 2'b01;
			14'b00101101100100: M1r = 2'b00;
			14'b01101101100100: M1r = 2'b00;
			14'b10101101100100: M1r = 2'b01;
			14'b11101101100100: M1r = 2'b01;
			14'b00111101100100: M1r = 2'b00;
			14'b01111101100100: M1r = 2'b00;
			14'b10111101100100: M1r = 2'b00;
			14'b11111101100100: M1r = 2'b00;
			14'b00000010100100: M1r = 2'b00;
			14'b01000010100100: M1r = 2'b00;
			14'b10000010100100: M1r = 2'b00;
			14'b11000010100100: M1r = 2'b00;
			14'b00010010100100: M1r = 2'b00;
			14'b01010010100100: M1r = 2'b00;
			14'b10010010100100: M1r = 2'b00;
			14'b11010010100100: M1r = 2'b00;
			14'b00100010100100: M1r = 2'b00;
			14'b01100010100100: M1r = 2'b00;
			14'b10100010100100: M1r = 2'b00;
			14'b11100010100100: M1r = 2'b00;
			14'b00110010100100: M1r = 2'b00;
			14'b01110010100100: M1r = 2'b00;
			14'b10110010100100: M1r = 2'b00;
			14'b11110010100100: M1r = 2'b00;
			14'b00000110100100: M1r = 2'b00;
			14'b01000110100100: M1r = 2'b00;
			14'b10000110100100: M1r = 2'b00;
			14'b11000110100100: M1r = 2'b00;
			14'b00010110100100: M1r = 2'b00;
			14'b01010110100100: M1r = 2'b00;
			14'b10010110100100: M1r = 2'b00;
			14'b11010110100100: M1r = 2'b00;
			14'b00100110100100: M1r = 2'b00;
			14'b01100110100100: M1r = 2'b00;
			14'b10100110100100: M1r = 2'b00;
			14'b11100110100100: M1r = 2'b00;
			14'b00110110100100: M1r = 2'b00;
			14'b01110110100100: M1r = 2'b00;
			14'b10110110100100: M1r = 2'b00;
			14'b11110110100100: M1r = 2'b00;
			14'b00001010100100: M1r = 2'b00;
			14'b01001010100100: M1r = 2'b00;
			14'b10001010100100: M1r = 2'b00;
			14'b11001010100100: M1r = 2'b01;
			14'b00011010100100: M1r = 2'b00;
			14'b01011010100100: M1r = 2'b00;
			14'b10011010100100: M1r = 2'b00;
			14'b11011010100100: M1r = 2'b00;
			14'b00101010100100: M1r = 2'b00;
			14'b01101010100100: M1r = 2'b00;
			14'b10101010100100: M1r = 2'b00;
			14'b11101010100100: M1r = 2'b00;
			14'b00111010100100: M1r = 2'b00;
			14'b01111010100100: M1r = 2'b00;
			14'b10111010100100: M1r = 2'b00;
			14'b11111010100100: M1r = 2'b00;
			14'b00001110100100: M1r = 2'b01;
			14'b01001110100100: M1r = 2'b01;
			14'b10001110100100: M1r = 2'b01;
			14'b11001110100100: M1r = 2'b01;
			14'b00011110100100: M1r = 2'b00;
			14'b01011110100100: M1r = 2'b01;
			14'b10011110100100: M1r = 2'b01;
			14'b11011110100100: M1r = 2'b01;
			14'b00101110100100: M1r = 2'b00;
			14'b01101110100100: M1r = 2'b00;
			14'b10101110100100: M1r = 2'b00;
			14'b11101110100100: M1r = 2'b00;
			14'b00111110100100: M1r = 2'b00;
			14'b01111110100100: M1r = 2'b00;
			14'b10111110100100: M1r = 2'b00;
			14'b11111110100100: M1r = 2'b00;
			14'b00000011100100: M1r = 2'b00;
			14'b01000011100100: M1r = 2'b00;
			14'b10000011100100: M1r = 2'b00;
			14'b11000011100100: M1r = 2'b00;
			14'b00010011100100: M1r = 2'b00;
			14'b01010011100100: M1r = 2'b00;
			14'b10010011100100: M1r = 2'b00;
			14'b11010011100100: M1r = 2'b00;
			14'b00100011100100: M1r = 2'b00;
			14'b01100011100100: M1r = 2'b00;
			14'b10100011100100: M1r = 2'b00;
			14'b11100011100100: M1r = 2'b00;
			14'b00110011100100: M1r = 2'b00;
			14'b01110011100100: M1r = 2'b00;
			14'b10110011100100: M1r = 2'b00;
			14'b11110011100100: M1r = 2'b00;
			14'b00000111100100: M1r = 2'b00;
			14'b01000111100100: M1r = 2'b00;
			14'b10000111100100: M1r = 2'b00;
			14'b11000111100100: M1r = 2'b00;
			14'b00010111100100: M1r = 2'b00;
			14'b01010111100100: M1r = 2'b00;
			14'b10010111100100: M1r = 2'b00;
			14'b11010111100100: M1r = 2'b00;
			14'b00100111100100: M1r = 2'b00;
			14'b01100111100100: M1r = 2'b00;
			14'b10100111100100: M1r = 2'b00;
			14'b11100111100100: M1r = 2'b00;
			14'b00110111100100: M1r = 2'b00;
			14'b01110111100100: M1r = 2'b00;
			14'b10110111100100: M1r = 2'b00;
			14'b11110111100100: M1r = 2'b00;
			14'b00001011100100: M1r = 2'b00;
			14'b01001011100100: M1r = 2'b00;
			14'b10001011100100: M1r = 2'b00;
			14'b11001011100100: M1r = 2'b00;
			14'b00011011100100: M1r = 2'b00;
			14'b01011011100100: M1r = 2'b00;
			14'b10011011100100: M1r = 2'b00;
			14'b11011011100100: M1r = 2'b00;
			14'b00101011100100: M1r = 2'b00;
			14'b01101011100100: M1r = 2'b00;
			14'b10101011100100: M1r = 2'b00;
			14'b11101011100100: M1r = 2'b00;
			14'b00111011100100: M1r = 2'b00;
			14'b01111011100100: M1r = 2'b00;
			14'b10111011100100: M1r = 2'b00;
			14'b11111011100100: M1r = 2'b00;
			14'b00001111100100: M1r = 2'b01;
			14'b01001111100100: M1r = 2'b01;
			14'b10001111100100: M1r = 2'b01;
			14'b11001111100100: M1r = 2'b01;
			14'b00011111100100: M1r = 2'b00;
			14'b01011111100100: M1r = 2'b00;
			14'b10011111100100: M1r = 2'b00;
			14'b11011111100100: M1r = 2'b01;
			14'b00101111100100: M1r = 2'b00;
			14'b01101111100100: M1r = 2'b00;
			14'b10101111100100: M1r = 2'b00;
			14'b11101111100100: M1r = 2'b00;
			14'b00111111100100: M1r = 2'b00;
			14'b01111111100100: M1r = 2'b00;
			14'b10111111100100: M1r = 2'b00;
			14'b11111111100100: M1r = 2'b00;
			14'b00000000110100: M1r = 2'b00;
			14'b01000000110100: M1r = 2'b00;
			14'b10000000110100: M1r = 2'b00;
			14'b11000000110100: M1r = 2'b00;
			14'b00010000110100: M1r = 2'b00;
			14'b01010000110100: M1r = 2'b00;
			14'b10010000110100: M1r = 2'b00;
			14'b11010000110100: M1r = 2'b00;
			14'b00100000110100: M1r = 2'b00;
			14'b01100000110100: M1r = 2'b00;
			14'b10100000110100: M1r = 2'b00;
			14'b11100000110100: M1r = 2'b00;
			14'b00110000110100: M1r = 2'b00;
			14'b01110000110100: M1r = 2'b00;
			14'b10110000110100: M1r = 2'b00;
			14'b11110000110100: M1r = 2'b00;
			14'b00000100110100: M1r = 2'b00;
			14'b01000100110100: M1r = 2'b01;
			14'b10000100110100: M1r = 2'b01;
			14'b11000100110100: M1r = 2'b01;
			14'b00010100110100: M1r = 2'b00;
			14'b01010100110100: M1r = 2'b00;
			14'b10010100110100: M1r = 2'b00;
			14'b11010100110100: M1r = 2'b00;
			14'b00100100110100: M1r = 2'b00;
			14'b01100100110100: M1r = 2'b00;
			14'b10100100110100: M1r = 2'b00;
			14'b11100100110100: M1r = 2'b00;
			14'b00110100110100: M1r = 2'b00;
			14'b01110100110100: M1r = 2'b00;
			14'b10110100110100: M1r = 2'b00;
			14'b11110100110100: M1r = 2'b00;
			14'b00001000110100: M1r = 2'b01;
			14'b01001000110100: M1r = 2'b01;
			14'b10001000110100: M1r = 2'b01;
			14'b11001000110100: M1r = 2'b10;
			14'b00011000110100: M1r = 2'b01;
			14'b01011000110100: M1r = 2'b01;
			14'b10011000110100: M1r = 2'b01;
			14'b11011000110100: M1r = 2'b01;
			14'b00101000110100: M1r = 2'b00;
			14'b01101000110100: M1r = 2'b00;
			14'b10101000110100: M1r = 2'b01;
			14'b11101000110100: M1r = 2'b01;
			14'b00111000110100: M1r = 2'b00;
			14'b01111000110100: M1r = 2'b00;
			14'b10111000110100: M1r = 2'b00;
			14'b11111000110100: M1r = 2'b00;
			14'b00001100110100: M1r = 2'b10;
			14'b01001100110100: M1r = 2'b10;
			14'b10001100110100: M1r = 2'b10;
			14'b11001100110100: M1r = 2'b10;
			14'b00011100110100: M1r = 2'b01;
			14'b01011100110100: M1r = 2'b10;
			14'b10011100110100: M1r = 2'b10;
			14'b11011100110100: M1r = 2'b10;
			14'b00101100110100: M1r = 2'b01;
			14'b01101100110100: M1r = 2'b01;
			14'b10101100110100: M1r = 2'b01;
			14'b11101100110100: M1r = 2'b01;
			14'b00111100110100: M1r = 2'b00;
			14'b01111100110100: M1r = 2'b01;
			14'b10111100110100: M1r = 2'b01;
			14'b11111100110100: M1r = 2'b01;
			14'b00000001110100: M1r = 2'b00;
			14'b01000001110100: M1r = 2'b00;
			14'b10000001110100: M1r = 2'b00;
			14'b11000001110100: M1r = 2'b00;
			14'b00010001110100: M1r = 2'b00;
			14'b01010001110100: M1r = 2'b00;
			14'b10010001110100: M1r = 2'b00;
			14'b11010001110100: M1r = 2'b00;
			14'b00100001110100: M1r = 2'b00;
			14'b01100001110100: M1r = 2'b00;
			14'b10100001110100: M1r = 2'b00;
			14'b11100001110100: M1r = 2'b00;
			14'b00110001110100: M1r = 2'b00;
			14'b01110001110100: M1r = 2'b00;
			14'b10110001110100: M1r = 2'b00;
			14'b11110001110100: M1r = 2'b00;
			14'b00000101110100: M1r = 2'b00;
			14'b01000101110100: M1r = 2'b00;
			14'b10000101110100: M1r = 2'b00;
			14'b11000101110100: M1r = 2'b01;
			14'b00010101110100: M1r = 2'b00;
			14'b01010101110100: M1r = 2'b00;
			14'b10010101110100: M1r = 2'b00;
			14'b11010101110100: M1r = 2'b00;
			14'b00100101110100: M1r = 2'b00;
			14'b01100101110100: M1r = 2'b00;
			14'b10100101110100: M1r = 2'b00;
			14'b11100101110100: M1r = 2'b00;
			14'b00110101110100: M1r = 2'b00;
			14'b01110101110100: M1r = 2'b00;
			14'b10110101110100: M1r = 2'b00;
			14'b11110101110100: M1r = 2'b00;
			14'b00001001110100: M1r = 2'b01;
			14'b01001001110100: M1r = 2'b01;
			14'b10001001110100: M1r = 2'b01;
			14'b11001001110100: M1r = 2'b01;
			14'b00011001110100: M1r = 2'b00;
			14'b01011001110100: M1r = 2'b01;
			14'b10011001110100: M1r = 2'b01;
			14'b11011001110100: M1r = 2'b01;
			14'b00101001110100: M1r = 2'b00;
			14'b01101001110100: M1r = 2'b00;
			14'b10101001110100: M1r = 2'b00;
			14'b11101001110100: M1r = 2'b00;
			14'b00111001110100: M1r = 2'b00;
			14'b01111001110100: M1r = 2'b00;
			14'b10111001110100: M1r = 2'b00;
			14'b11111001110100: M1r = 2'b00;
			14'b00001101110100: M1r = 2'b10;
			14'b01001101110100: M1r = 2'b10;
			14'b10001101110100: M1r = 2'b10;
			14'b11001101110100: M1r = 2'b10;
			14'b00011101110100: M1r = 2'b01;
			14'b01011101110100: M1r = 2'b01;
			14'b10011101110100: M1r = 2'b01;
			14'b11011101110100: M1r = 2'b10;
			14'b00101101110100: M1r = 2'b01;
			14'b01101101110100: M1r = 2'b01;
			14'b10101101110100: M1r = 2'b01;
			14'b11101101110100: M1r = 2'b01;
			14'b00111101110100: M1r = 2'b00;
			14'b01111101110100: M1r = 2'b00;
			14'b10111101110100: M1r = 2'b01;
			14'b11111101110100: M1r = 2'b01;
			14'b00000010110100: M1r = 2'b00;
			14'b01000010110100: M1r = 2'b00;
			14'b10000010110100: M1r = 2'b00;
			14'b11000010110100: M1r = 2'b00;
			14'b00010010110100: M1r = 2'b00;
			14'b01010010110100: M1r = 2'b00;
			14'b10010010110100: M1r = 2'b00;
			14'b11010010110100: M1r = 2'b00;
			14'b00100010110100: M1r = 2'b00;
			14'b01100010110100: M1r = 2'b00;
			14'b10100010110100: M1r = 2'b00;
			14'b11100010110100: M1r = 2'b00;
			14'b00110010110100: M1r = 2'b00;
			14'b01110010110100: M1r = 2'b00;
			14'b10110010110100: M1r = 2'b00;
			14'b11110010110100: M1r = 2'b00;
			14'b00000110110100: M1r = 2'b00;
			14'b01000110110100: M1r = 2'b00;
			14'b10000110110100: M1r = 2'b00;
			14'b11000110110100: M1r = 2'b00;
			14'b00010110110100: M1r = 2'b00;
			14'b01010110110100: M1r = 2'b00;
			14'b10010110110100: M1r = 2'b00;
			14'b11010110110100: M1r = 2'b00;
			14'b00100110110100: M1r = 2'b00;
			14'b01100110110100: M1r = 2'b00;
			14'b10100110110100: M1r = 2'b00;
			14'b11100110110100: M1r = 2'b00;
			14'b00110110110100: M1r = 2'b00;
			14'b01110110110100: M1r = 2'b00;
			14'b10110110110100: M1r = 2'b00;
			14'b11110110110100: M1r = 2'b00;
			14'b00001010110100: M1r = 2'b01;
			14'b01001010110100: M1r = 2'b01;
			14'b10001010110100: M1r = 2'b01;
			14'b11001010110100: M1r = 2'b01;
			14'b00011010110100: M1r = 2'b00;
			14'b01011010110100: M1r = 2'b00;
			14'b10011010110100: M1r = 2'b00;
			14'b11011010110100: M1r = 2'b01;
			14'b00101010110100: M1r = 2'b00;
			14'b01101010110100: M1r = 2'b00;
			14'b10101010110100: M1r = 2'b00;
			14'b11101010110100: M1r = 2'b00;
			14'b00111010110100: M1r = 2'b00;
			14'b01111010110100: M1r = 2'b00;
			14'b10111010110100: M1r = 2'b00;
			14'b11111010110100: M1r = 2'b00;
			14'b00001110110100: M1r = 2'b01;
			14'b01001110110100: M1r = 2'b10;
			14'b10001110110100: M1r = 2'b10;
			14'b11001110110100: M1r = 2'b10;
			14'b00011110110100: M1r = 2'b01;
			14'b01011110110100: M1r = 2'b01;
			14'b10011110110100: M1r = 2'b01;
			14'b11011110110100: M1r = 2'b01;
			14'b00101110110100: M1r = 2'b00;
			14'b01101110110100: M1r = 2'b01;
			14'b10101110110100: M1r = 2'b01;
			14'b11101110110100: M1r = 2'b01;
			14'b00111110110100: M1r = 2'b00;
			14'b01111110110100: M1r = 2'b00;
			14'b10111110110100: M1r = 2'b00;
			14'b11111110110100: M1r = 2'b00;
			14'b00000011110100: M1r = 2'b00;
			14'b01000011110100: M1r = 2'b00;
			14'b10000011110100: M1r = 2'b00;
			14'b11000011110100: M1r = 2'b00;
			14'b00010011110100: M1r = 2'b00;
			14'b01010011110100: M1r = 2'b00;
			14'b10010011110100: M1r = 2'b00;
			14'b11010011110100: M1r = 2'b00;
			14'b00100011110100: M1r = 2'b00;
			14'b01100011110100: M1r = 2'b00;
			14'b10100011110100: M1r = 2'b00;
			14'b11100011110100: M1r = 2'b00;
			14'b00110011110100: M1r = 2'b00;
			14'b01110011110100: M1r = 2'b00;
			14'b10110011110100: M1r = 2'b00;
			14'b11110011110100: M1r = 2'b00;
			14'b00000111110100: M1r = 2'b00;
			14'b01000111110100: M1r = 2'b00;
			14'b10000111110100: M1r = 2'b00;
			14'b11000111110100: M1r = 2'b00;
			14'b00010111110100: M1r = 2'b00;
			14'b01010111110100: M1r = 2'b00;
			14'b10010111110100: M1r = 2'b00;
			14'b11010111110100: M1r = 2'b00;
			14'b00100111110100: M1r = 2'b00;
			14'b01100111110100: M1r = 2'b00;
			14'b10100111110100: M1r = 2'b00;
			14'b11100111110100: M1r = 2'b00;
			14'b00110111110100: M1r = 2'b00;
			14'b01110111110100: M1r = 2'b00;
			14'b10110111110100: M1r = 2'b00;
			14'b11110111110100: M1r = 2'b00;
			14'b00001011110100: M1r = 2'b00;
			14'b01001011110100: M1r = 2'b00;
			14'b10001011110100: M1r = 2'b01;
			14'b11001011110100: M1r = 2'b01;
			14'b00011011110100: M1r = 2'b00;
			14'b01011011110100: M1r = 2'b00;
			14'b10011011110100: M1r = 2'b00;
			14'b11011011110100: M1r = 2'b00;
			14'b00101011110100: M1r = 2'b00;
			14'b01101011110100: M1r = 2'b00;
			14'b10101011110100: M1r = 2'b00;
			14'b11101011110100: M1r = 2'b00;
			14'b00111011110100: M1r = 2'b00;
			14'b01111011110100: M1r = 2'b00;
			14'b10111011110100: M1r = 2'b00;
			14'b11111011110100: M1r = 2'b00;
			14'b00001111110100: M1r = 2'b01;
			14'b01001111110100: M1r = 2'b01;
			14'b10001111110100: M1r = 2'b01;
			14'b11001111110100: M1r = 2'b10;
			14'b00011111110100: M1r = 2'b01;
			14'b01011111110100: M1r = 2'b01;
			14'b10011111110100: M1r = 2'b01;
			14'b11011111110100: M1r = 2'b01;
			14'b00101111110100: M1r = 2'b00;
			14'b01101111110100: M1r = 2'b00;
			14'b10101111110100: M1r = 2'b00;
			14'b11101111110100: M1r = 2'b01;
			14'b00111111110100: M1r = 2'b00;
			14'b01111111110100: M1r = 2'b00;
			14'b10111111110100: M1r = 2'b00;
			14'b11111111110100: M1r = 2'b00;
			14'b00000000001000: M1r = 2'b00;
			14'b01000000001000: M1r = 2'b00;
			14'b10000000001000: M1r = 2'b00;
			14'b11000000001000: M1r = 2'b00;
			14'b00010000001000: M1r = 2'b00;
			14'b01010000001000: M1r = 2'b00;
			14'b10010000001000: M1r = 2'b00;
			14'b11010000001000: M1r = 2'b00;
			14'b00100000001000: M1r = 2'b00;
			14'b01100000001000: M1r = 2'b00;
			14'b10100000001000: M1r = 2'b00;
			14'b11100000001000: M1r = 2'b00;
			14'b00110000001000: M1r = 2'b00;
			14'b01110000001000: M1r = 2'b00;
			14'b10110000001000: M1r = 2'b00;
			14'b11110000001000: M1r = 2'b00;
			14'b00000100001000: M1r = 2'b00;
			14'b01000100001000: M1r = 2'b00;
			14'b10000100001000: M1r = 2'b00;
			14'b11000100001000: M1r = 2'b00;
			14'b00010100001000: M1r = 2'b00;
			14'b01010100001000: M1r = 2'b00;
			14'b10010100001000: M1r = 2'b00;
			14'b11010100001000: M1r = 2'b00;
			14'b00100100001000: M1r = 2'b00;
			14'b01100100001000: M1r = 2'b00;
			14'b10100100001000: M1r = 2'b00;
			14'b11100100001000: M1r = 2'b00;
			14'b00110100001000: M1r = 2'b00;
			14'b01110100001000: M1r = 2'b00;
			14'b10110100001000: M1r = 2'b00;
			14'b11110100001000: M1r = 2'b00;
			14'b00001000001000: M1r = 2'b00;
			14'b01001000001000: M1r = 2'b00;
			14'b10001000001000: M1r = 2'b00;
			14'b11001000001000: M1r = 2'b00;
			14'b00011000001000: M1r = 2'b00;
			14'b01011000001000: M1r = 2'b00;
			14'b10011000001000: M1r = 2'b00;
			14'b11011000001000: M1r = 2'b00;
			14'b00101000001000: M1r = 2'b00;
			14'b01101000001000: M1r = 2'b00;
			14'b10101000001000: M1r = 2'b00;
			14'b11101000001000: M1r = 2'b00;
			14'b00111000001000: M1r = 2'b00;
			14'b01111000001000: M1r = 2'b00;
			14'b10111000001000: M1r = 2'b00;
			14'b11111000001000: M1r = 2'b00;
			14'b00001100001000: M1r = 2'b00;
			14'b01001100001000: M1r = 2'b00;
			14'b10001100001000: M1r = 2'b00;
			14'b11001100001000: M1r = 2'b00;
			14'b00011100001000: M1r = 2'b00;
			14'b01011100001000: M1r = 2'b00;
			14'b10011100001000: M1r = 2'b00;
			14'b11011100001000: M1r = 2'b00;
			14'b00101100001000: M1r = 2'b00;
			14'b01101100001000: M1r = 2'b00;
			14'b10101100001000: M1r = 2'b00;
			14'b11101100001000: M1r = 2'b00;
			14'b00111100001000: M1r = 2'b00;
			14'b01111100001000: M1r = 2'b00;
			14'b10111100001000: M1r = 2'b00;
			14'b11111100001000: M1r = 2'b00;
			14'b00000001001000: M1r = 2'b00;
			14'b01000001001000: M1r = 2'b00;
			14'b10000001001000: M1r = 2'b00;
			14'b11000001001000: M1r = 2'b00;
			14'b00010001001000: M1r = 2'b00;
			14'b01010001001000: M1r = 2'b00;
			14'b10010001001000: M1r = 2'b00;
			14'b11010001001000: M1r = 2'b00;
			14'b00100001001000: M1r = 2'b00;
			14'b01100001001000: M1r = 2'b00;
			14'b10100001001000: M1r = 2'b00;
			14'b11100001001000: M1r = 2'b00;
			14'b00110001001000: M1r = 2'b00;
			14'b01110001001000: M1r = 2'b00;
			14'b10110001001000: M1r = 2'b00;
			14'b11110001001000: M1r = 2'b00;
			14'b00000101001000: M1r = 2'b00;
			14'b01000101001000: M1r = 2'b00;
			14'b10000101001000: M1r = 2'b00;
			14'b11000101001000: M1r = 2'b00;
			14'b00010101001000: M1r = 2'b00;
			14'b01010101001000: M1r = 2'b00;
			14'b10010101001000: M1r = 2'b00;
			14'b11010101001000: M1r = 2'b00;
			14'b00100101001000: M1r = 2'b00;
			14'b01100101001000: M1r = 2'b00;
			14'b10100101001000: M1r = 2'b00;
			14'b11100101001000: M1r = 2'b00;
			14'b00110101001000: M1r = 2'b00;
			14'b01110101001000: M1r = 2'b00;
			14'b10110101001000: M1r = 2'b00;
			14'b11110101001000: M1r = 2'b00;
			14'b00001001001000: M1r = 2'b00;
			14'b01001001001000: M1r = 2'b00;
			14'b10001001001000: M1r = 2'b00;
			14'b11001001001000: M1r = 2'b00;
			14'b00011001001000: M1r = 2'b00;
			14'b01011001001000: M1r = 2'b00;
			14'b10011001001000: M1r = 2'b00;
			14'b11011001001000: M1r = 2'b00;
			14'b00101001001000: M1r = 2'b00;
			14'b01101001001000: M1r = 2'b00;
			14'b10101001001000: M1r = 2'b00;
			14'b11101001001000: M1r = 2'b00;
			14'b00111001001000: M1r = 2'b00;
			14'b01111001001000: M1r = 2'b00;
			14'b10111001001000: M1r = 2'b00;
			14'b11111001001000: M1r = 2'b00;
			14'b00001101001000: M1r = 2'b00;
			14'b01001101001000: M1r = 2'b00;
			14'b10001101001000: M1r = 2'b00;
			14'b11001101001000: M1r = 2'b00;
			14'b00011101001000: M1r = 2'b00;
			14'b01011101001000: M1r = 2'b00;
			14'b10011101001000: M1r = 2'b00;
			14'b11011101001000: M1r = 2'b00;
			14'b00101101001000: M1r = 2'b00;
			14'b01101101001000: M1r = 2'b00;
			14'b10101101001000: M1r = 2'b00;
			14'b11101101001000: M1r = 2'b00;
			14'b00111101001000: M1r = 2'b00;
			14'b01111101001000: M1r = 2'b00;
			14'b10111101001000: M1r = 2'b00;
			14'b11111101001000: M1r = 2'b00;
			14'b00000010001000: M1r = 2'b00;
			14'b01000010001000: M1r = 2'b00;
			14'b10000010001000: M1r = 2'b00;
			14'b11000010001000: M1r = 2'b00;
			14'b00010010001000: M1r = 2'b00;
			14'b01010010001000: M1r = 2'b00;
			14'b10010010001000: M1r = 2'b00;
			14'b11010010001000: M1r = 2'b00;
			14'b00100010001000: M1r = 2'b00;
			14'b01100010001000: M1r = 2'b00;
			14'b10100010001000: M1r = 2'b00;
			14'b11100010001000: M1r = 2'b00;
			14'b00110010001000: M1r = 2'b00;
			14'b01110010001000: M1r = 2'b00;
			14'b10110010001000: M1r = 2'b00;
			14'b11110010001000: M1r = 2'b00;
			14'b00000110001000: M1r = 2'b00;
			14'b01000110001000: M1r = 2'b00;
			14'b10000110001000: M1r = 2'b00;
			14'b11000110001000: M1r = 2'b00;
			14'b00010110001000: M1r = 2'b00;
			14'b01010110001000: M1r = 2'b00;
			14'b10010110001000: M1r = 2'b00;
			14'b11010110001000: M1r = 2'b00;
			14'b00100110001000: M1r = 2'b00;
			14'b01100110001000: M1r = 2'b00;
			14'b10100110001000: M1r = 2'b00;
			14'b11100110001000: M1r = 2'b00;
			14'b00110110001000: M1r = 2'b00;
			14'b01110110001000: M1r = 2'b00;
			14'b10110110001000: M1r = 2'b00;
			14'b11110110001000: M1r = 2'b00;
			14'b00001010001000: M1r = 2'b00;
			14'b01001010001000: M1r = 2'b00;
			14'b10001010001000: M1r = 2'b00;
			14'b11001010001000: M1r = 2'b00;
			14'b00011010001000: M1r = 2'b00;
			14'b01011010001000: M1r = 2'b00;
			14'b10011010001000: M1r = 2'b00;
			14'b11011010001000: M1r = 2'b00;
			14'b00101010001000: M1r = 2'b00;
			14'b01101010001000: M1r = 2'b00;
			14'b10101010001000: M1r = 2'b00;
			14'b11101010001000: M1r = 2'b00;
			14'b00111010001000: M1r = 2'b00;
			14'b01111010001000: M1r = 2'b00;
			14'b10111010001000: M1r = 2'b00;
			14'b11111010001000: M1r = 2'b00;
			14'b00001110001000: M1r = 2'b00;
			14'b01001110001000: M1r = 2'b00;
			14'b10001110001000: M1r = 2'b00;
			14'b11001110001000: M1r = 2'b00;
			14'b00011110001000: M1r = 2'b00;
			14'b01011110001000: M1r = 2'b00;
			14'b10011110001000: M1r = 2'b00;
			14'b11011110001000: M1r = 2'b00;
			14'b00101110001000: M1r = 2'b00;
			14'b01101110001000: M1r = 2'b00;
			14'b10101110001000: M1r = 2'b00;
			14'b11101110001000: M1r = 2'b00;
			14'b00111110001000: M1r = 2'b00;
			14'b01111110001000: M1r = 2'b00;
			14'b10111110001000: M1r = 2'b00;
			14'b11111110001000: M1r = 2'b00;
			14'b00000011001000: M1r = 2'b00;
			14'b01000011001000: M1r = 2'b00;
			14'b10000011001000: M1r = 2'b00;
			14'b11000011001000: M1r = 2'b00;
			14'b00010011001000: M1r = 2'b00;
			14'b01010011001000: M1r = 2'b00;
			14'b10010011001000: M1r = 2'b00;
			14'b11010011001000: M1r = 2'b00;
			14'b00100011001000: M1r = 2'b00;
			14'b01100011001000: M1r = 2'b00;
			14'b10100011001000: M1r = 2'b00;
			14'b11100011001000: M1r = 2'b00;
			14'b00110011001000: M1r = 2'b00;
			14'b01110011001000: M1r = 2'b00;
			14'b10110011001000: M1r = 2'b00;
			14'b11110011001000: M1r = 2'b00;
			14'b00000111001000: M1r = 2'b00;
			14'b01000111001000: M1r = 2'b00;
			14'b10000111001000: M1r = 2'b00;
			14'b11000111001000: M1r = 2'b00;
			14'b00010111001000: M1r = 2'b00;
			14'b01010111001000: M1r = 2'b00;
			14'b10010111001000: M1r = 2'b00;
			14'b11010111001000: M1r = 2'b00;
			14'b00100111001000: M1r = 2'b00;
			14'b01100111001000: M1r = 2'b00;
			14'b10100111001000: M1r = 2'b00;
			14'b11100111001000: M1r = 2'b00;
			14'b00110111001000: M1r = 2'b00;
			14'b01110111001000: M1r = 2'b00;
			14'b10110111001000: M1r = 2'b00;
			14'b11110111001000: M1r = 2'b00;
			14'b00001011001000: M1r = 2'b00;
			14'b01001011001000: M1r = 2'b00;
			14'b10001011001000: M1r = 2'b00;
			14'b11001011001000: M1r = 2'b00;
			14'b00011011001000: M1r = 2'b00;
			14'b01011011001000: M1r = 2'b00;
			14'b10011011001000: M1r = 2'b00;
			14'b11011011001000: M1r = 2'b00;
			14'b00101011001000: M1r = 2'b00;
			14'b01101011001000: M1r = 2'b00;
			14'b10101011001000: M1r = 2'b00;
			14'b11101011001000: M1r = 2'b00;
			14'b00111011001000: M1r = 2'b00;
			14'b01111011001000: M1r = 2'b00;
			14'b10111011001000: M1r = 2'b00;
			14'b11111011001000: M1r = 2'b00;
			14'b00001111001000: M1r = 2'b00;
			14'b01001111001000: M1r = 2'b00;
			14'b10001111001000: M1r = 2'b00;
			14'b11001111001000: M1r = 2'b00;
			14'b00011111001000: M1r = 2'b00;
			14'b01011111001000: M1r = 2'b00;
			14'b10011111001000: M1r = 2'b00;
			14'b11011111001000: M1r = 2'b00;
			14'b00101111001000: M1r = 2'b00;
			14'b01101111001000: M1r = 2'b00;
			14'b10101111001000: M1r = 2'b00;
			14'b11101111001000: M1r = 2'b00;
			14'b00111111001000: M1r = 2'b00;
			14'b01111111001000: M1r = 2'b00;
			14'b10111111001000: M1r = 2'b00;
			14'b11111111001000: M1r = 2'b00;
			14'b00000000011000: M1r = 2'b00;
			14'b01000000011000: M1r = 2'b00;
			14'b10000000011000: M1r = 2'b00;
			14'b11000000011000: M1r = 2'b00;
			14'b00010000011000: M1r = 2'b00;
			14'b01010000011000: M1r = 2'b00;
			14'b10010000011000: M1r = 2'b00;
			14'b11010000011000: M1r = 2'b00;
			14'b00100000011000: M1r = 2'b00;
			14'b01100000011000: M1r = 2'b00;
			14'b10100000011000: M1r = 2'b00;
			14'b11100000011000: M1r = 2'b00;
			14'b00110000011000: M1r = 2'b00;
			14'b01110000011000: M1r = 2'b00;
			14'b10110000011000: M1r = 2'b00;
			14'b11110000011000: M1r = 2'b00;
			14'b00000100011000: M1r = 2'b00;
			14'b01000100011000: M1r = 2'b00;
			14'b10000100011000: M1r = 2'b00;
			14'b11000100011000: M1r = 2'b00;
			14'b00010100011000: M1r = 2'b00;
			14'b01010100011000: M1r = 2'b00;
			14'b10010100011000: M1r = 2'b00;
			14'b11010100011000: M1r = 2'b00;
			14'b00100100011000: M1r = 2'b00;
			14'b01100100011000: M1r = 2'b00;
			14'b10100100011000: M1r = 2'b00;
			14'b11100100011000: M1r = 2'b00;
			14'b00110100011000: M1r = 2'b00;
			14'b01110100011000: M1r = 2'b00;
			14'b10110100011000: M1r = 2'b00;
			14'b11110100011000: M1r = 2'b00;
			14'b00001000011000: M1r = 2'b00;
			14'b01001000011000: M1r = 2'b00;
			14'b10001000011000: M1r = 2'b00;
			14'b11001000011000: M1r = 2'b00;
			14'b00011000011000: M1r = 2'b00;
			14'b01011000011000: M1r = 2'b00;
			14'b10011000011000: M1r = 2'b00;
			14'b11011000011000: M1r = 2'b00;
			14'b00101000011000: M1r = 2'b00;
			14'b01101000011000: M1r = 2'b00;
			14'b10101000011000: M1r = 2'b00;
			14'b11101000011000: M1r = 2'b00;
			14'b00111000011000: M1r = 2'b00;
			14'b01111000011000: M1r = 2'b00;
			14'b10111000011000: M1r = 2'b00;
			14'b11111000011000: M1r = 2'b00;
			14'b00001100011000: M1r = 2'b00;
			14'b01001100011000: M1r = 2'b00;
			14'b10001100011000: M1r = 2'b01;
			14'b11001100011000: M1r = 2'b01;
			14'b00011100011000: M1r = 2'b00;
			14'b01011100011000: M1r = 2'b00;
			14'b10011100011000: M1r = 2'b00;
			14'b11011100011000: M1r = 2'b00;
			14'b00101100011000: M1r = 2'b00;
			14'b01101100011000: M1r = 2'b00;
			14'b10101100011000: M1r = 2'b00;
			14'b11101100011000: M1r = 2'b00;
			14'b00111100011000: M1r = 2'b00;
			14'b01111100011000: M1r = 2'b00;
			14'b10111100011000: M1r = 2'b00;
			14'b11111100011000: M1r = 2'b00;
			14'b00000001011000: M1r = 2'b00;
			14'b01000001011000: M1r = 2'b00;
			14'b10000001011000: M1r = 2'b00;
			14'b11000001011000: M1r = 2'b00;
			14'b00010001011000: M1r = 2'b00;
			14'b01010001011000: M1r = 2'b00;
			14'b10010001011000: M1r = 2'b00;
			14'b11010001011000: M1r = 2'b00;
			14'b00100001011000: M1r = 2'b00;
			14'b01100001011000: M1r = 2'b00;
			14'b10100001011000: M1r = 2'b00;
			14'b11100001011000: M1r = 2'b00;
			14'b00110001011000: M1r = 2'b00;
			14'b01110001011000: M1r = 2'b00;
			14'b10110001011000: M1r = 2'b00;
			14'b11110001011000: M1r = 2'b00;
			14'b00000101011000: M1r = 2'b00;
			14'b01000101011000: M1r = 2'b00;
			14'b10000101011000: M1r = 2'b00;
			14'b11000101011000: M1r = 2'b00;
			14'b00010101011000: M1r = 2'b00;
			14'b01010101011000: M1r = 2'b00;
			14'b10010101011000: M1r = 2'b00;
			14'b11010101011000: M1r = 2'b00;
			14'b00100101011000: M1r = 2'b00;
			14'b01100101011000: M1r = 2'b00;
			14'b10100101011000: M1r = 2'b00;
			14'b11100101011000: M1r = 2'b00;
			14'b00110101011000: M1r = 2'b00;
			14'b01110101011000: M1r = 2'b00;
			14'b10110101011000: M1r = 2'b00;
			14'b11110101011000: M1r = 2'b00;
			14'b00001001011000: M1r = 2'b00;
			14'b01001001011000: M1r = 2'b00;
			14'b10001001011000: M1r = 2'b00;
			14'b11001001011000: M1r = 2'b00;
			14'b00011001011000: M1r = 2'b00;
			14'b01011001011000: M1r = 2'b00;
			14'b10011001011000: M1r = 2'b00;
			14'b11011001011000: M1r = 2'b00;
			14'b00101001011000: M1r = 2'b00;
			14'b01101001011000: M1r = 2'b00;
			14'b10101001011000: M1r = 2'b00;
			14'b11101001011000: M1r = 2'b00;
			14'b00111001011000: M1r = 2'b00;
			14'b01111001011000: M1r = 2'b00;
			14'b10111001011000: M1r = 2'b00;
			14'b11111001011000: M1r = 2'b00;
			14'b00001101011000: M1r = 2'b00;
			14'b01001101011000: M1r = 2'b00;
			14'b10001101011000: M1r = 2'b00;
			14'b11001101011000: M1r = 2'b00;
			14'b00011101011000: M1r = 2'b00;
			14'b01011101011000: M1r = 2'b00;
			14'b10011101011000: M1r = 2'b00;
			14'b11011101011000: M1r = 2'b00;
			14'b00101101011000: M1r = 2'b00;
			14'b01101101011000: M1r = 2'b00;
			14'b10101101011000: M1r = 2'b00;
			14'b11101101011000: M1r = 2'b00;
			14'b00111101011000: M1r = 2'b00;
			14'b01111101011000: M1r = 2'b00;
			14'b10111101011000: M1r = 2'b00;
			14'b11111101011000: M1r = 2'b00;
			14'b00000010011000: M1r = 2'b00;
			14'b01000010011000: M1r = 2'b00;
			14'b10000010011000: M1r = 2'b00;
			14'b11000010011000: M1r = 2'b00;
			14'b00010010011000: M1r = 2'b00;
			14'b01010010011000: M1r = 2'b00;
			14'b10010010011000: M1r = 2'b00;
			14'b11010010011000: M1r = 2'b00;
			14'b00100010011000: M1r = 2'b00;
			14'b01100010011000: M1r = 2'b00;
			14'b10100010011000: M1r = 2'b00;
			14'b11100010011000: M1r = 2'b00;
			14'b00110010011000: M1r = 2'b00;
			14'b01110010011000: M1r = 2'b00;
			14'b10110010011000: M1r = 2'b00;
			14'b11110010011000: M1r = 2'b00;
			14'b00000110011000: M1r = 2'b00;
			14'b01000110011000: M1r = 2'b00;
			14'b10000110011000: M1r = 2'b00;
			14'b11000110011000: M1r = 2'b00;
			14'b00010110011000: M1r = 2'b00;
			14'b01010110011000: M1r = 2'b00;
			14'b10010110011000: M1r = 2'b00;
			14'b11010110011000: M1r = 2'b00;
			14'b00100110011000: M1r = 2'b00;
			14'b01100110011000: M1r = 2'b00;
			14'b10100110011000: M1r = 2'b00;
			14'b11100110011000: M1r = 2'b00;
			14'b00110110011000: M1r = 2'b00;
			14'b01110110011000: M1r = 2'b00;
			14'b10110110011000: M1r = 2'b00;
			14'b11110110011000: M1r = 2'b00;
			14'b00001010011000: M1r = 2'b00;
			14'b01001010011000: M1r = 2'b00;
			14'b10001010011000: M1r = 2'b00;
			14'b11001010011000: M1r = 2'b00;
			14'b00011010011000: M1r = 2'b00;
			14'b01011010011000: M1r = 2'b00;
			14'b10011010011000: M1r = 2'b00;
			14'b11011010011000: M1r = 2'b00;
			14'b00101010011000: M1r = 2'b00;
			14'b01101010011000: M1r = 2'b00;
			14'b10101010011000: M1r = 2'b00;
			14'b11101010011000: M1r = 2'b00;
			14'b00111010011000: M1r = 2'b00;
			14'b01111010011000: M1r = 2'b00;
			14'b10111010011000: M1r = 2'b00;
			14'b11111010011000: M1r = 2'b00;
			14'b00001110011000: M1r = 2'b00;
			14'b01001110011000: M1r = 2'b00;
			14'b10001110011000: M1r = 2'b00;
			14'b11001110011000: M1r = 2'b00;
			14'b00011110011000: M1r = 2'b00;
			14'b01011110011000: M1r = 2'b00;
			14'b10011110011000: M1r = 2'b00;
			14'b11011110011000: M1r = 2'b00;
			14'b00101110011000: M1r = 2'b00;
			14'b01101110011000: M1r = 2'b00;
			14'b10101110011000: M1r = 2'b00;
			14'b11101110011000: M1r = 2'b00;
			14'b00111110011000: M1r = 2'b00;
			14'b01111110011000: M1r = 2'b00;
			14'b10111110011000: M1r = 2'b00;
			14'b11111110011000: M1r = 2'b00;
			14'b00000011011000: M1r = 2'b00;
			14'b01000011011000: M1r = 2'b00;
			14'b10000011011000: M1r = 2'b00;
			14'b11000011011000: M1r = 2'b00;
			14'b00010011011000: M1r = 2'b00;
			14'b01010011011000: M1r = 2'b00;
			14'b10010011011000: M1r = 2'b00;
			14'b11010011011000: M1r = 2'b00;
			14'b00100011011000: M1r = 2'b00;
			14'b01100011011000: M1r = 2'b00;
			14'b10100011011000: M1r = 2'b00;
			14'b11100011011000: M1r = 2'b00;
			14'b00110011011000: M1r = 2'b00;
			14'b01110011011000: M1r = 2'b00;
			14'b10110011011000: M1r = 2'b00;
			14'b11110011011000: M1r = 2'b00;
			14'b00000111011000: M1r = 2'b00;
			14'b01000111011000: M1r = 2'b00;
			14'b10000111011000: M1r = 2'b00;
			14'b11000111011000: M1r = 2'b00;
			14'b00010111011000: M1r = 2'b00;
			14'b01010111011000: M1r = 2'b00;
			14'b10010111011000: M1r = 2'b00;
			14'b11010111011000: M1r = 2'b00;
			14'b00100111011000: M1r = 2'b00;
			14'b01100111011000: M1r = 2'b00;
			14'b10100111011000: M1r = 2'b00;
			14'b11100111011000: M1r = 2'b00;
			14'b00110111011000: M1r = 2'b00;
			14'b01110111011000: M1r = 2'b00;
			14'b10110111011000: M1r = 2'b00;
			14'b11110111011000: M1r = 2'b00;
			14'b00001011011000: M1r = 2'b00;
			14'b01001011011000: M1r = 2'b00;
			14'b10001011011000: M1r = 2'b00;
			14'b11001011011000: M1r = 2'b00;
			14'b00011011011000: M1r = 2'b00;
			14'b01011011011000: M1r = 2'b00;
			14'b10011011011000: M1r = 2'b00;
			14'b11011011011000: M1r = 2'b00;
			14'b00101011011000: M1r = 2'b00;
			14'b01101011011000: M1r = 2'b00;
			14'b10101011011000: M1r = 2'b00;
			14'b11101011011000: M1r = 2'b00;
			14'b00111011011000: M1r = 2'b00;
			14'b01111011011000: M1r = 2'b00;
			14'b10111011011000: M1r = 2'b00;
			14'b11111011011000: M1r = 2'b00;
			14'b00001111011000: M1r = 2'b00;
			14'b01001111011000: M1r = 2'b00;
			14'b10001111011000: M1r = 2'b00;
			14'b11001111011000: M1r = 2'b00;
			14'b00011111011000: M1r = 2'b00;
			14'b01011111011000: M1r = 2'b00;
			14'b10011111011000: M1r = 2'b00;
			14'b11011111011000: M1r = 2'b00;
			14'b00101111011000: M1r = 2'b00;
			14'b01101111011000: M1r = 2'b00;
			14'b10101111011000: M1r = 2'b00;
			14'b11101111011000: M1r = 2'b00;
			14'b00111111011000: M1r = 2'b00;
			14'b01111111011000: M1r = 2'b00;
			14'b10111111011000: M1r = 2'b00;
			14'b11111111011000: M1r = 2'b00;
			14'b00000000101000: M1r = 2'b00;
			14'b01000000101000: M1r = 2'b00;
			14'b10000000101000: M1r = 2'b00;
			14'b11000000101000: M1r = 2'b00;
			14'b00010000101000: M1r = 2'b00;
			14'b01010000101000: M1r = 2'b00;
			14'b10010000101000: M1r = 2'b00;
			14'b11010000101000: M1r = 2'b00;
			14'b00100000101000: M1r = 2'b00;
			14'b01100000101000: M1r = 2'b00;
			14'b10100000101000: M1r = 2'b00;
			14'b11100000101000: M1r = 2'b00;
			14'b00110000101000: M1r = 2'b00;
			14'b01110000101000: M1r = 2'b00;
			14'b10110000101000: M1r = 2'b00;
			14'b11110000101000: M1r = 2'b00;
			14'b00000100101000: M1r = 2'b00;
			14'b01000100101000: M1r = 2'b00;
			14'b10000100101000: M1r = 2'b00;
			14'b11000100101000: M1r = 2'b00;
			14'b00010100101000: M1r = 2'b00;
			14'b01010100101000: M1r = 2'b00;
			14'b10010100101000: M1r = 2'b00;
			14'b11010100101000: M1r = 2'b00;
			14'b00100100101000: M1r = 2'b00;
			14'b01100100101000: M1r = 2'b00;
			14'b10100100101000: M1r = 2'b00;
			14'b11100100101000: M1r = 2'b00;
			14'b00110100101000: M1r = 2'b00;
			14'b01110100101000: M1r = 2'b00;
			14'b10110100101000: M1r = 2'b00;
			14'b11110100101000: M1r = 2'b00;
			14'b00001000101000: M1r = 2'b00;
			14'b01001000101000: M1r = 2'b00;
			14'b10001000101000: M1r = 2'b00;
			14'b11001000101000: M1r = 2'b00;
			14'b00011000101000: M1r = 2'b00;
			14'b01011000101000: M1r = 2'b00;
			14'b10011000101000: M1r = 2'b00;
			14'b11011000101000: M1r = 2'b00;
			14'b00101000101000: M1r = 2'b00;
			14'b01101000101000: M1r = 2'b00;
			14'b10101000101000: M1r = 2'b00;
			14'b11101000101000: M1r = 2'b00;
			14'b00111000101000: M1r = 2'b00;
			14'b01111000101000: M1r = 2'b00;
			14'b10111000101000: M1r = 2'b00;
			14'b11111000101000: M1r = 2'b00;
			14'b00001100101000: M1r = 2'b01;
			14'b01001100101000: M1r = 2'b01;
			14'b10001100101000: M1r = 2'b01;
			14'b11001100101000: M1r = 2'b01;
			14'b00011100101000: M1r = 2'b00;
			14'b01011100101000: M1r = 2'b00;
			14'b10011100101000: M1r = 2'b01;
			14'b11011100101000: M1r = 2'b01;
			14'b00101100101000: M1r = 2'b00;
			14'b01101100101000: M1r = 2'b00;
			14'b10101100101000: M1r = 2'b00;
			14'b11101100101000: M1r = 2'b00;
			14'b00111100101000: M1r = 2'b00;
			14'b01111100101000: M1r = 2'b00;
			14'b10111100101000: M1r = 2'b00;
			14'b11111100101000: M1r = 2'b00;
			14'b00000001101000: M1r = 2'b00;
			14'b01000001101000: M1r = 2'b00;
			14'b10000001101000: M1r = 2'b00;
			14'b11000001101000: M1r = 2'b00;
			14'b00010001101000: M1r = 2'b00;
			14'b01010001101000: M1r = 2'b00;
			14'b10010001101000: M1r = 2'b00;
			14'b11010001101000: M1r = 2'b00;
			14'b00100001101000: M1r = 2'b00;
			14'b01100001101000: M1r = 2'b00;
			14'b10100001101000: M1r = 2'b00;
			14'b11100001101000: M1r = 2'b00;
			14'b00110001101000: M1r = 2'b00;
			14'b01110001101000: M1r = 2'b00;
			14'b10110001101000: M1r = 2'b00;
			14'b11110001101000: M1r = 2'b00;
			14'b00000101101000: M1r = 2'b00;
			14'b01000101101000: M1r = 2'b00;
			14'b10000101101000: M1r = 2'b00;
			14'b11000101101000: M1r = 2'b00;
			14'b00010101101000: M1r = 2'b00;
			14'b01010101101000: M1r = 2'b00;
			14'b10010101101000: M1r = 2'b00;
			14'b11010101101000: M1r = 2'b00;
			14'b00100101101000: M1r = 2'b00;
			14'b01100101101000: M1r = 2'b00;
			14'b10100101101000: M1r = 2'b00;
			14'b11100101101000: M1r = 2'b00;
			14'b00110101101000: M1r = 2'b00;
			14'b01110101101000: M1r = 2'b00;
			14'b10110101101000: M1r = 2'b00;
			14'b11110101101000: M1r = 2'b00;
			14'b00001001101000: M1r = 2'b00;
			14'b01001001101000: M1r = 2'b00;
			14'b10001001101000: M1r = 2'b00;
			14'b11001001101000: M1r = 2'b00;
			14'b00011001101000: M1r = 2'b00;
			14'b01011001101000: M1r = 2'b00;
			14'b10011001101000: M1r = 2'b00;
			14'b11011001101000: M1r = 2'b00;
			14'b00101001101000: M1r = 2'b00;
			14'b01101001101000: M1r = 2'b00;
			14'b10101001101000: M1r = 2'b00;
			14'b11101001101000: M1r = 2'b00;
			14'b00111001101000: M1r = 2'b00;
			14'b01111001101000: M1r = 2'b00;
			14'b10111001101000: M1r = 2'b00;
			14'b11111001101000: M1r = 2'b00;
			14'b00001101101000: M1r = 2'b00;
			14'b01001101101000: M1r = 2'b01;
			14'b10001101101000: M1r = 2'b01;
			14'b11001101101000: M1r = 2'b01;
			14'b00011101101000: M1r = 2'b00;
			14'b01011101101000: M1r = 2'b00;
			14'b10011101101000: M1r = 2'b00;
			14'b11011101101000: M1r = 2'b00;
			14'b00101101101000: M1r = 2'b00;
			14'b01101101101000: M1r = 2'b00;
			14'b10101101101000: M1r = 2'b00;
			14'b11101101101000: M1r = 2'b00;
			14'b00111101101000: M1r = 2'b00;
			14'b01111101101000: M1r = 2'b00;
			14'b10111101101000: M1r = 2'b00;
			14'b11111101101000: M1r = 2'b00;
			14'b00000010101000: M1r = 2'b00;
			14'b01000010101000: M1r = 2'b00;
			14'b10000010101000: M1r = 2'b00;
			14'b11000010101000: M1r = 2'b00;
			14'b00010010101000: M1r = 2'b00;
			14'b01010010101000: M1r = 2'b00;
			14'b10010010101000: M1r = 2'b00;
			14'b11010010101000: M1r = 2'b00;
			14'b00100010101000: M1r = 2'b00;
			14'b01100010101000: M1r = 2'b00;
			14'b10100010101000: M1r = 2'b00;
			14'b11100010101000: M1r = 2'b00;
			14'b00110010101000: M1r = 2'b00;
			14'b01110010101000: M1r = 2'b00;
			14'b10110010101000: M1r = 2'b00;
			14'b11110010101000: M1r = 2'b00;
			14'b00000110101000: M1r = 2'b00;
			14'b01000110101000: M1r = 2'b00;
			14'b10000110101000: M1r = 2'b00;
			14'b11000110101000: M1r = 2'b00;
			14'b00010110101000: M1r = 2'b00;
			14'b01010110101000: M1r = 2'b00;
			14'b10010110101000: M1r = 2'b00;
			14'b11010110101000: M1r = 2'b00;
			14'b00100110101000: M1r = 2'b00;
			14'b01100110101000: M1r = 2'b00;
			14'b10100110101000: M1r = 2'b00;
			14'b11100110101000: M1r = 2'b00;
			14'b00110110101000: M1r = 2'b00;
			14'b01110110101000: M1r = 2'b00;
			14'b10110110101000: M1r = 2'b00;
			14'b11110110101000: M1r = 2'b00;
			14'b00001010101000: M1r = 2'b00;
			14'b01001010101000: M1r = 2'b00;
			14'b10001010101000: M1r = 2'b00;
			14'b11001010101000: M1r = 2'b00;
			14'b00011010101000: M1r = 2'b00;
			14'b01011010101000: M1r = 2'b00;
			14'b10011010101000: M1r = 2'b00;
			14'b11011010101000: M1r = 2'b00;
			14'b00101010101000: M1r = 2'b00;
			14'b01101010101000: M1r = 2'b00;
			14'b10101010101000: M1r = 2'b00;
			14'b11101010101000: M1r = 2'b00;
			14'b00111010101000: M1r = 2'b00;
			14'b01111010101000: M1r = 2'b00;
			14'b10111010101000: M1r = 2'b00;
			14'b11111010101000: M1r = 2'b00;
			14'b00001110101000: M1r = 2'b00;
			14'b01001110101000: M1r = 2'b00;
			14'b10001110101000: M1r = 2'b00;
			14'b11001110101000: M1r = 2'b01;
			14'b00011110101000: M1r = 2'b00;
			14'b01011110101000: M1r = 2'b00;
			14'b10011110101000: M1r = 2'b00;
			14'b11011110101000: M1r = 2'b00;
			14'b00101110101000: M1r = 2'b00;
			14'b01101110101000: M1r = 2'b00;
			14'b10101110101000: M1r = 2'b00;
			14'b11101110101000: M1r = 2'b00;
			14'b00111110101000: M1r = 2'b00;
			14'b01111110101000: M1r = 2'b00;
			14'b10111110101000: M1r = 2'b00;
			14'b11111110101000: M1r = 2'b00;
			14'b00000011101000: M1r = 2'b00;
			14'b01000011101000: M1r = 2'b00;
			14'b10000011101000: M1r = 2'b00;
			14'b11000011101000: M1r = 2'b00;
			14'b00010011101000: M1r = 2'b00;
			14'b01010011101000: M1r = 2'b00;
			14'b10010011101000: M1r = 2'b00;
			14'b11010011101000: M1r = 2'b00;
			14'b00100011101000: M1r = 2'b00;
			14'b01100011101000: M1r = 2'b00;
			14'b10100011101000: M1r = 2'b00;
			14'b11100011101000: M1r = 2'b00;
			14'b00110011101000: M1r = 2'b00;
			14'b01110011101000: M1r = 2'b00;
			14'b10110011101000: M1r = 2'b00;
			14'b11110011101000: M1r = 2'b00;
			14'b00000111101000: M1r = 2'b00;
			14'b01000111101000: M1r = 2'b00;
			14'b10000111101000: M1r = 2'b00;
			14'b11000111101000: M1r = 2'b00;
			14'b00010111101000: M1r = 2'b00;
			14'b01010111101000: M1r = 2'b00;
			14'b10010111101000: M1r = 2'b00;
			14'b11010111101000: M1r = 2'b00;
			14'b00100111101000: M1r = 2'b00;
			14'b01100111101000: M1r = 2'b00;
			14'b10100111101000: M1r = 2'b00;
			14'b11100111101000: M1r = 2'b00;
			14'b00110111101000: M1r = 2'b00;
			14'b01110111101000: M1r = 2'b00;
			14'b10110111101000: M1r = 2'b00;
			14'b11110111101000: M1r = 2'b00;
			14'b00001011101000: M1r = 2'b00;
			14'b01001011101000: M1r = 2'b00;
			14'b10001011101000: M1r = 2'b00;
			14'b11001011101000: M1r = 2'b00;
			14'b00011011101000: M1r = 2'b00;
			14'b01011011101000: M1r = 2'b00;
			14'b10011011101000: M1r = 2'b00;
			14'b11011011101000: M1r = 2'b00;
			14'b00101011101000: M1r = 2'b00;
			14'b01101011101000: M1r = 2'b00;
			14'b10101011101000: M1r = 2'b00;
			14'b11101011101000: M1r = 2'b00;
			14'b00111011101000: M1r = 2'b00;
			14'b01111011101000: M1r = 2'b00;
			14'b10111011101000: M1r = 2'b00;
			14'b11111011101000: M1r = 2'b00;
			14'b00001111101000: M1r = 2'b00;
			14'b01001111101000: M1r = 2'b00;
			14'b10001111101000: M1r = 2'b00;
			14'b11001111101000: M1r = 2'b00;
			14'b00011111101000: M1r = 2'b00;
			14'b01011111101000: M1r = 2'b00;
			14'b10011111101000: M1r = 2'b00;
			14'b11011111101000: M1r = 2'b00;
			14'b00101111101000: M1r = 2'b00;
			14'b01101111101000: M1r = 2'b00;
			14'b10101111101000: M1r = 2'b00;
			14'b11101111101000: M1r = 2'b00;
			14'b00111111101000: M1r = 2'b00;
			14'b01111111101000: M1r = 2'b00;
			14'b10111111101000: M1r = 2'b00;
			14'b11111111101000: M1r = 2'b00;
			14'b00000000111000: M1r = 2'b00;
			14'b01000000111000: M1r = 2'b00;
			14'b10000000111000: M1r = 2'b00;
			14'b11000000111000: M1r = 2'b00;
			14'b00010000111000: M1r = 2'b00;
			14'b01010000111000: M1r = 2'b00;
			14'b10010000111000: M1r = 2'b00;
			14'b11010000111000: M1r = 2'b00;
			14'b00100000111000: M1r = 2'b00;
			14'b01100000111000: M1r = 2'b00;
			14'b10100000111000: M1r = 2'b00;
			14'b11100000111000: M1r = 2'b00;
			14'b00110000111000: M1r = 2'b00;
			14'b01110000111000: M1r = 2'b00;
			14'b10110000111000: M1r = 2'b00;
			14'b11110000111000: M1r = 2'b00;
			14'b00000100111000: M1r = 2'b00;
			14'b01000100111000: M1r = 2'b00;
			14'b10000100111000: M1r = 2'b00;
			14'b11000100111000: M1r = 2'b00;
			14'b00010100111000: M1r = 2'b00;
			14'b01010100111000: M1r = 2'b00;
			14'b10010100111000: M1r = 2'b00;
			14'b11010100111000: M1r = 2'b00;
			14'b00100100111000: M1r = 2'b00;
			14'b01100100111000: M1r = 2'b00;
			14'b10100100111000: M1r = 2'b00;
			14'b11100100111000: M1r = 2'b00;
			14'b00110100111000: M1r = 2'b00;
			14'b01110100111000: M1r = 2'b00;
			14'b10110100111000: M1r = 2'b00;
			14'b11110100111000: M1r = 2'b00;
			14'b00001000111000: M1r = 2'b00;
			14'b01001000111000: M1r = 2'b01;
			14'b10001000111000: M1r = 2'b01;
			14'b11001000111000: M1r = 2'b01;
			14'b00011000111000: M1r = 2'b00;
			14'b01011000111000: M1r = 2'b00;
			14'b10011000111000: M1r = 2'b00;
			14'b11011000111000: M1r = 2'b00;
			14'b00101000111000: M1r = 2'b00;
			14'b01101000111000: M1r = 2'b00;
			14'b10101000111000: M1r = 2'b00;
			14'b11101000111000: M1r = 2'b00;
			14'b00111000111000: M1r = 2'b00;
			14'b01111000111000: M1r = 2'b00;
			14'b10111000111000: M1r = 2'b00;
			14'b11111000111000: M1r = 2'b00;
			14'b00001100111000: M1r = 2'b01;
			14'b01001100111000: M1r = 2'b01;
			14'b10001100111000: M1r = 2'b01;
			14'b11001100111000: M1r = 2'b10;
			14'b00011100111000: M1r = 2'b01;
			14'b01011100111000: M1r = 2'b01;
			14'b10011100111000: M1r = 2'b01;
			14'b11011100111000: M1r = 2'b01;
			14'b00101100111000: M1r = 2'b00;
			14'b01101100111000: M1r = 2'b00;
			14'b10101100111000: M1r = 2'b00;
			14'b11101100111000: M1r = 2'b01;
			14'b00111100111000: M1r = 2'b00;
			14'b01111100111000: M1r = 2'b00;
			14'b10111100111000: M1r = 2'b00;
			14'b11111100111000: M1r = 2'b00;
			14'b00000001111000: M1r = 2'b00;
			14'b01000001111000: M1r = 2'b00;
			14'b10000001111000: M1r = 2'b00;
			14'b11000001111000: M1r = 2'b00;
			14'b00010001111000: M1r = 2'b00;
			14'b01010001111000: M1r = 2'b00;
			14'b10010001111000: M1r = 2'b00;
			14'b11010001111000: M1r = 2'b00;
			14'b00100001111000: M1r = 2'b00;
			14'b01100001111000: M1r = 2'b00;
			14'b10100001111000: M1r = 2'b00;
			14'b11100001111000: M1r = 2'b00;
			14'b00110001111000: M1r = 2'b00;
			14'b01110001111000: M1r = 2'b00;
			14'b10110001111000: M1r = 2'b00;
			14'b11110001111000: M1r = 2'b00;
			14'b00000101111000: M1r = 2'b00;
			14'b01000101111000: M1r = 2'b00;
			14'b10000101111000: M1r = 2'b00;
			14'b11000101111000: M1r = 2'b00;
			14'b00010101111000: M1r = 2'b00;
			14'b01010101111000: M1r = 2'b00;
			14'b10010101111000: M1r = 2'b00;
			14'b11010101111000: M1r = 2'b00;
			14'b00100101111000: M1r = 2'b00;
			14'b01100101111000: M1r = 2'b00;
			14'b10100101111000: M1r = 2'b00;
			14'b11100101111000: M1r = 2'b00;
			14'b00110101111000: M1r = 2'b00;
			14'b01110101111000: M1r = 2'b00;
			14'b10110101111000: M1r = 2'b00;
			14'b11110101111000: M1r = 2'b00;
			14'b00001001111000: M1r = 2'b00;
			14'b01001001111000: M1r = 2'b00;
			14'b10001001111000: M1r = 2'b00;
			14'b11001001111000: M1r = 2'b01;
			14'b00011001111000: M1r = 2'b00;
			14'b01011001111000: M1r = 2'b00;
			14'b10011001111000: M1r = 2'b00;
			14'b11011001111000: M1r = 2'b00;
			14'b00101001111000: M1r = 2'b00;
			14'b01101001111000: M1r = 2'b00;
			14'b10101001111000: M1r = 2'b00;
			14'b11101001111000: M1r = 2'b00;
			14'b00111001111000: M1r = 2'b00;
			14'b01111001111000: M1r = 2'b00;
			14'b10111001111000: M1r = 2'b00;
			14'b11111001111000: M1r = 2'b00;
			14'b00001101111000: M1r = 2'b01;
			14'b01001101111000: M1r = 2'b01;
			14'b10001101111000: M1r = 2'b01;
			14'b11001101111000: M1r = 2'b01;
			14'b00011101111000: M1r = 2'b00;
			14'b01011101111000: M1r = 2'b01;
			14'b10011101111000: M1r = 2'b01;
			14'b11011101111000: M1r = 2'b01;
			14'b00101101111000: M1r = 2'b00;
			14'b01101101111000: M1r = 2'b00;
			14'b10101101111000: M1r = 2'b00;
			14'b11101101111000: M1r = 2'b00;
			14'b00111101111000: M1r = 2'b00;
			14'b01111101111000: M1r = 2'b00;
			14'b10111101111000: M1r = 2'b00;
			14'b11111101111000: M1r = 2'b00;
			14'b00000010111000: M1r = 2'b00;
			14'b01000010111000: M1r = 2'b00;
			14'b10000010111000: M1r = 2'b00;
			14'b11000010111000: M1r = 2'b00;
			14'b00010010111000: M1r = 2'b00;
			14'b01010010111000: M1r = 2'b00;
			14'b10010010111000: M1r = 2'b00;
			14'b11010010111000: M1r = 2'b00;
			14'b00100010111000: M1r = 2'b00;
			14'b01100010111000: M1r = 2'b00;
			14'b10100010111000: M1r = 2'b00;
			14'b11100010111000: M1r = 2'b00;
			14'b00110010111000: M1r = 2'b00;
			14'b01110010111000: M1r = 2'b00;
			14'b10110010111000: M1r = 2'b00;
			14'b11110010111000: M1r = 2'b00;
			14'b00000110111000: M1r = 2'b00;
			14'b01000110111000: M1r = 2'b00;
			14'b10000110111000: M1r = 2'b00;
			14'b11000110111000: M1r = 2'b00;
			14'b00010110111000: M1r = 2'b00;
			14'b01010110111000: M1r = 2'b00;
			14'b10010110111000: M1r = 2'b00;
			14'b11010110111000: M1r = 2'b00;
			14'b00100110111000: M1r = 2'b00;
			14'b01100110111000: M1r = 2'b00;
			14'b10100110111000: M1r = 2'b00;
			14'b11100110111000: M1r = 2'b00;
			14'b00110110111000: M1r = 2'b00;
			14'b01110110111000: M1r = 2'b00;
			14'b10110110111000: M1r = 2'b00;
			14'b11110110111000: M1r = 2'b00;
			14'b00001010111000: M1r = 2'b00;
			14'b01001010111000: M1r = 2'b00;
			14'b10001010111000: M1r = 2'b00;
			14'b11001010111000: M1r = 2'b00;
			14'b00011010111000: M1r = 2'b00;
			14'b01011010111000: M1r = 2'b00;
			14'b10011010111000: M1r = 2'b00;
			14'b11011010111000: M1r = 2'b00;
			14'b00101010111000: M1r = 2'b00;
			14'b01101010111000: M1r = 2'b00;
			14'b10101010111000: M1r = 2'b00;
			14'b11101010111000: M1r = 2'b00;
			14'b00111010111000: M1r = 2'b00;
			14'b01111010111000: M1r = 2'b00;
			14'b10111010111000: M1r = 2'b00;
			14'b11111010111000: M1r = 2'b00;
			14'b00001110111000: M1r = 2'b01;
			14'b01001110111000: M1r = 2'b01;
			14'b10001110111000: M1r = 2'b01;
			14'b11001110111000: M1r = 2'b01;
			14'b00011110111000: M1r = 2'b00;
			14'b01011110111000: M1r = 2'b00;
			14'b10011110111000: M1r = 2'b00;
			14'b11011110111000: M1r = 2'b01;
			14'b00101110111000: M1r = 2'b00;
			14'b01101110111000: M1r = 2'b00;
			14'b10101110111000: M1r = 2'b00;
			14'b11101110111000: M1r = 2'b00;
			14'b00111110111000: M1r = 2'b00;
			14'b01111110111000: M1r = 2'b00;
			14'b10111110111000: M1r = 2'b00;
			14'b11111110111000: M1r = 2'b00;
			14'b00000011111000: M1r = 2'b00;
			14'b01000011111000: M1r = 2'b00;
			14'b10000011111000: M1r = 2'b00;
			14'b11000011111000: M1r = 2'b00;
			14'b00010011111000: M1r = 2'b00;
			14'b01010011111000: M1r = 2'b00;
			14'b10010011111000: M1r = 2'b00;
			14'b11010011111000: M1r = 2'b00;
			14'b00100011111000: M1r = 2'b00;
			14'b01100011111000: M1r = 2'b00;
			14'b10100011111000: M1r = 2'b00;
			14'b11100011111000: M1r = 2'b00;
			14'b00110011111000: M1r = 2'b00;
			14'b01110011111000: M1r = 2'b00;
			14'b10110011111000: M1r = 2'b00;
			14'b11110011111000: M1r = 2'b00;
			14'b00000111111000: M1r = 2'b00;
			14'b01000111111000: M1r = 2'b00;
			14'b10000111111000: M1r = 2'b00;
			14'b11000111111000: M1r = 2'b00;
			14'b00010111111000: M1r = 2'b00;
			14'b01010111111000: M1r = 2'b00;
			14'b10010111111000: M1r = 2'b00;
			14'b11010111111000: M1r = 2'b00;
			14'b00100111111000: M1r = 2'b00;
			14'b01100111111000: M1r = 2'b00;
			14'b10100111111000: M1r = 2'b00;
			14'b11100111111000: M1r = 2'b00;
			14'b00110111111000: M1r = 2'b00;
			14'b01110111111000: M1r = 2'b00;
			14'b10110111111000: M1r = 2'b00;
			14'b11110111111000: M1r = 2'b00;
			14'b00001011111000: M1r = 2'b00;
			14'b01001011111000: M1r = 2'b00;
			14'b10001011111000: M1r = 2'b00;
			14'b11001011111000: M1r = 2'b00;
			14'b00011011111000: M1r = 2'b00;
			14'b01011011111000: M1r = 2'b00;
			14'b10011011111000: M1r = 2'b00;
			14'b11011011111000: M1r = 2'b00;
			14'b00101011111000: M1r = 2'b00;
			14'b01101011111000: M1r = 2'b00;
			14'b10101011111000: M1r = 2'b00;
			14'b11101011111000: M1r = 2'b00;
			14'b00111011111000: M1r = 2'b00;
			14'b01111011111000: M1r = 2'b00;
			14'b10111011111000: M1r = 2'b00;
			14'b11111011111000: M1r = 2'b00;
			14'b00001111111000: M1r = 2'b00;
			14'b01001111111000: M1r = 2'b00;
			14'b10001111111000: M1r = 2'b01;
			14'b11001111111000: M1r = 2'b01;
			14'b00011111111000: M1r = 2'b00;
			14'b01011111111000: M1r = 2'b00;
			14'b10011111111000: M1r = 2'b00;
			14'b11011111111000: M1r = 2'b00;
			14'b00101111111000: M1r = 2'b00;
			14'b01101111111000: M1r = 2'b00;
			14'b10101111111000: M1r = 2'b00;
			14'b11101111111000: M1r = 2'b00;
			14'b00111111111000: M1r = 2'b00;
			14'b01111111111000: M1r = 2'b00;
			14'b10111111111000: M1r = 2'b00;
			14'b11111111111000: M1r = 2'b00;
			14'b00000000001100: M1r = 2'b00;
			14'b01000000001100: M1r = 2'b00;
			14'b10000000001100: M1r = 2'b00;
			14'b11000000001100: M1r = 2'b00;
			14'b00010000001100: M1r = 2'b00;
			14'b01010000001100: M1r = 2'b00;
			14'b10010000001100: M1r = 2'b00;
			14'b11010000001100: M1r = 2'b00;
			14'b00100000001100: M1r = 2'b00;
			14'b01100000001100: M1r = 2'b00;
			14'b10100000001100: M1r = 2'b00;
			14'b11100000001100: M1r = 2'b00;
			14'b00110000001100: M1r = 2'b00;
			14'b01110000001100: M1r = 2'b00;
			14'b10110000001100: M1r = 2'b00;
			14'b11110000001100: M1r = 2'b00;
			14'b00000100001100: M1r = 2'b00;
			14'b01000100001100: M1r = 2'b00;
			14'b10000100001100: M1r = 2'b00;
			14'b11000100001100: M1r = 2'b00;
			14'b00010100001100: M1r = 2'b00;
			14'b01010100001100: M1r = 2'b00;
			14'b10010100001100: M1r = 2'b00;
			14'b11010100001100: M1r = 2'b00;
			14'b00100100001100: M1r = 2'b00;
			14'b01100100001100: M1r = 2'b00;
			14'b10100100001100: M1r = 2'b00;
			14'b11100100001100: M1r = 2'b00;
			14'b00110100001100: M1r = 2'b00;
			14'b01110100001100: M1r = 2'b00;
			14'b10110100001100: M1r = 2'b00;
			14'b11110100001100: M1r = 2'b00;
			14'b00001000001100: M1r = 2'b00;
			14'b01001000001100: M1r = 2'b00;
			14'b10001000001100: M1r = 2'b00;
			14'b11001000001100: M1r = 2'b00;
			14'b00011000001100: M1r = 2'b00;
			14'b01011000001100: M1r = 2'b00;
			14'b10011000001100: M1r = 2'b00;
			14'b11011000001100: M1r = 2'b00;
			14'b00101000001100: M1r = 2'b00;
			14'b01101000001100: M1r = 2'b00;
			14'b10101000001100: M1r = 2'b00;
			14'b11101000001100: M1r = 2'b00;
			14'b00111000001100: M1r = 2'b00;
			14'b01111000001100: M1r = 2'b00;
			14'b10111000001100: M1r = 2'b00;
			14'b11111000001100: M1r = 2'b00;
			14'b00001100001100: M1r = 2'b00;
			14'b01001100001100: M1r = 2'b00;
			14'b10001100001100: M1r = 2'b00;
			14'b11001100001100: M1r = 2'b00;
			14'b00011100001100: M1r = 2'b00;
			14'b01011100001100: M1r = 2'b00;
			14'b10011100001100: M1r = 2'b00;
			14'b11011100001100: M1r = 2'b00;
			14'b00101100001100: M1r = 2'b00;
			14'b01101100001100: M1r = 2'b00;
			14'b10101100001100: M1r = 2'b00;
			14'b11101100001100: M1r = 2'b00;
			14'b00111100001100: M1r = 2'b00;
			14'b01111100001100: M1r = 2'b00;
			14'b10111100001100: M1r = 2'b00;
			14'b11111100001100: M1r = 2'b00;
			14'b00000001001100: M1r = 2'b00;
			14'b01000001001100: M1r = 2'b00;
			14'b10000001001100: M1r = 2'b00;
			14'b11000001001100: M1r = 2'b00;
			14'b00010001001100: M1r = 2'b00;
			14'b01010001001100: M1r = 2'b00;
			14'b10010001001100: M1r = 2'b00;
			14'b11010001001100: M1r = 2'b00;
			14'b00100001001100: M1r = 2'b00;
			14'b01100001001100: M1r = 2'b00;
			14'b10100001001100: M1r = 2'b00;
			14'b11100001001100: M1r = 2'b00;
			14'b00110001001100: M1r = 2'b00;
			14'b01110001001100: M1r = 2'b00;
			14'b10110001001100: M1r = 2'b00;
			14'b11110001001100: M1r = 2'b00;
			14'b00000101001100: M1r = 2'b00;
			14'b01000101001100: M1r = 2'b00;
			14'b10000101001100: M1r = 2'b00;
			14'b11000101001100: M1r = 2'b00;
			14'b00010101001100: M1r = 2'b00;
			14'b01010101001100: M1r = 2'b00;
			14'b10010101001100: M1r = 2'b00;
			14'b11010101001100: M1r = 2'b00;
			14'b00100101001100: M1r = 2'b00;
			14'b01100101001100: M1r = 2'b00;
			14'b10100101001100: M1r = 2'b00;
			14'b11100101001100: M1r = 2'b00;
			14'b00110101001100: M1r = 2'b00;
			14'b01110101001100: M1r = 2'b00;
			14'b10110101001100: M1r = 2'b00;
			14'b11110101001100: M1r = 2'b00;
			14'b00001001001100: M1r = 2'b00;
			14'b01001001001100: M1r = 2'b00;
			14'b10001001001100: M1r = 2'b00;
			14'b11001001001100: M1r = 2'b00;
			14'b00011001001100: M1r = 2'b00;
			14'b01011001001100: M1r = 2'b00;
			14'b10011001001100: M1r = 2'b00;
			14'b11011001001100: M1r = 2'b00;
			14'b00101001001100: M1r = 2'b00;
			14'b01101001001100: M1r = 2'b00;
			14'b10101001001100: M1r = 2'b00;
			14'b11101001001100: M1r = 2'b00;
			14'b00111001001100: M1r = 2'b00;
			14'b01111001001100: M1r = 2'b00;
			14'b10111001001100: M1r = 2'b00;
			14'b11111001001100: M1r = 2'b00;
			14'b00001101001100: M1r = 2'b00;
			14'b01001101001100: M1r = 2'b00;
			14'b10001101001100: M1r = 2'b00;
			14'b11001101001100: M1r = 2'b00;
			14'b00011101001100: M1r = 2'b00;
			14'b01011101001100: M1r = 2'b00;
			14'b10011101001100: M1r = 2'b00;
			14'b11011101001100: M1r = 2'b00;
			14'b00101101001100: M1r = 2'b00;
			14'b01101101001100: M1r = 2'b00;
			14'b10101101001100: M1r = 2'b00;
			14'b11101101001100: M1r = 2'b00;
			14'b00111101001100: M1r = 2'b00;
			14'b01111101001100: M1r = 2'b00;
			14'b10111101001100: M1r = 2'b00;
			14'b11111101001100: M1r = 2'b00;
			14'b00000010001100: M1r = 2'b00;
			14'b01000010001100: M1r = 2'b00;
			14'b10000010001100: M1r = 2'b00;
			14'b11000010001100: M1r = 2'b00;
			14'b00010010001100: M1r = 2'b00;
			14'b01010010001100: M1r = 2'b00;
			14'b10010010001100: M1r = 2'b00;
			14'b11010010001100: M1r = 2'b00;
			14'b00100010001100: M1r = 2'b00;
			14'b01100010001100: M1r = 2'b00;
			14'b10100010001100: M1r = 2'b00;
			14'b11100010001100: M1r = 2'b00;
			14'b00110010001100: M1r = 2'b00;
			14'b01110010001100: M1r = 2'b00;
			14'b10110010001100: M1r = 2'b00;
			14'b11110010001100: M1r = 2'b00;
			14'b00000110001100: M1r = 2'b00;
			14'b01000110001100: M1r = 2'b00;
			14'b10000110001100: M1r = 2'b00;
			14'b11000110001100: M1r = 2'b00;
			14'b00010110001100: M1r = 2'b00;
			14'b01010110001100: M1r = 2'b00;
			14'b10010110001100: M1r = 2'b00;
			14'b11010110001100: M1r = 2'b00;
			14'b00100110001100: M1r = 2'b00;
			14'b01100110001100: M1r = 2'b00;
			14'b10100110001100: M1r = 2'b00;
			14'b11100110001100: M1r = 2'b00;
			14'b00110110001100: M1r = 2'b00;
			14'b01110110001100: M1r = 2'b00;
			14'b10110110001100: M1r = 2'b00;
			14'b11110110001100: M1r = 2'b00;
			14'b00001010001100: M1r = 2'b00;
			14'b01001010001100: M1r = 2'b00;
			14'b10001010001100: M1r = 2'b00;
			14'b11001010001100: M1r = 2'b00;
			14'b00011010001100: M1r = 2'b00;
			14'b01011010001100: M1r = 2'b00;
			14'b10011010001100: M1r = 2'b00;
			14'b11011010001100: M1r = 2'b00;
			14'b00101010001100: M1r = 2'b00;
			14'b01101010001100: M1r = 2'b00;
			14'b10101010001100: M1r = 2'b00;
			14'b11101010001100: M1r = 2'b00;
			14'b00111010001100: M1r = 2'b00;
			14'b01111010001100: M1r = 2'b00;
			14'b10111010001100: M1r = 2'b00;
			14'b11111010001100: M1r = 2'b00;
			14'b00001110001100: M1r = 2'b00;
			14'b01001110001100: M1r = 2'b00;
			14'b10001110001100: M1r = 2'b00;
			14'b11001110001100: M1r = 2'b00;
			14'b00011110001100: M1r = 2'b00;
			14'b01011110001100: M1r = 2'b00;
			14'b10011110001100: M1r = 2'b00;
			14'b11011110001100: M1r = 2'b00;
			14'b00101110001100: M1r = 2'b00;
			14'b01101110001100: M1r = 2'b00;
			14'b10101110001100: M1r = 2'b00;
			14'b11101110001100: M1r = 2'b00;
			14'b00111110001100: M1r = 2'b00;
			14'b01111110001100: M1r = 2'b00;
			14'b10111110001100: M1r = 2'b00;
			14'b11111110001100: M1r = 2'b00;
			14'b00000011001100: M1r = 2'b00;
			14'b01000011001100: M1r = 2'b00;
			14'b10000011001100: M1r = 2'b00;
			14'b11000011001100: M1r = 2'b00;
			14'b00010011001100: M1r = 2'b00;
			14'b01010011001100: M1r = 2'b00;
			14'b10010011001100: M1r = 2'b00;
			14'b11010011001100: M1r = 2'b00;
			14'b00100011001100: M1r = 2'b00;
			14'b01100011001100: M1r = 2'b00;
			14'b10100011001100: M1r = 2'b00;
			14'b11100011001100: M1r = 2'b00;
			14'b00110011001100: M1r = 2'b00;
			14'b01110011001100: M1r = 2'b00;
			14'b10110011001100: M1r = 2'b00;
			14'b11110011001100: M1r = 2'b00;
			14'b00000111001100: M1r = 2'b00;
			14'b01000111001100: M1r = 2'b00;
			14'b10000111001100: M1r = 2'b00;
			14'b11000111001100: M1r = 2'b00;
			14'b00010111001100: M1r = 2'b00;
			14'b01010111001100: M1r = 2'b00;
			14'b10010111001100: M1r = 2'b00;
			14'b11010111001100: M1r = 2'b00;
			14'b00100111001100: M1r = 2'b00;
			14'b01100111001100: M1r = 2'b00;
			14'b10100111001100: M1r = 2'b00;
			14'b11100111001100: M1r = 2'b00;
			14'b00110111001100: M1r = 2'b00;
			14'b01110111001100: M1r = 2'b00;
			14'b10110111001100: M1r = 2'b00;
			14'b11110111001100: M1r = 2'b00;
			14'b00001011001100: M1r = 2'b00;
			14'b01001011001100: M1r = 2'b00;
			14'b10001011001100: M1r = 2'b00;
			14'b11001011001100: M1r = 2'b00;
			14'b00011011001100: M1r = 2'b00;
			14'b01011011001100: M1r = 2'b00;
			14'b10011011001100: M1r = 2'b00;
			14'b11011011001100: M1r = 2'b00;
			14'b00101011001100: M1r = 2'b00;
			14'b01101011001100: M1r = 2'b00;
			14'b10101011001100: M1r = 2'b00;
			14'b11101011001100: M1r = 2'b00;
			14'b00111011001100: M1r = 2'b00;
			14'b01111011001100: M1r = 2'b00;
			14'b10111011001100: M1r = 2'b00;
			14'b11111011001100: M1r = 2'b00;
			14'b00001111001100: M1r = 2'b00;
			14'b01001111001100: M1r = 2'b00;
			14'b10001111001100: M1r = 2'b00;
			14'b11001111001100: M1r = 2'b00;
			14'b00011111001100: M1r = 2'b00;
			14'b01011111001100: M1r = 2'b00;
			14'b10011111001100: M1r = 2'b00;
			14'b11011111001100: M1r = 2'b00;
			14'b00101111001100: M1r = 2'b00;
			14'b01101111001100: M1r = 2'b00;
			14'b10101111001100: M1r = 2'b00;
			14'b11101111001100: M1r = 2'b00;
			14'b00111111001100: M1r = 2'b00;
			14'b01111111001100: M1r = 2'b00;
			14'b10111111001100: M1r = 2'b00;
			14'b11111111001100: M1r = 2'b00;
			14'b00000000011100: M1r = 2'b00;
			14'b01000000011100: M1r = 2'b00;
			14'b10000000011100: M1r = 2'b00;
			14'b11000000011100: M1r = 2'b00;
			14'b00010000011100: M1r = 2'b00;
			14'b01010000011100: M1r = 2'b00;
			14'b10010000011100: M1r = 2'b00;
			14'b11010000011100: M1r = 2'b00;
			14'b00100000011100: M1r = 2'b00;
			14'b01100000011100: M1r = 2'b00;
			14'b10100000011100: M1r = 2'b00;
			14'b11100000011100: M1r = 2'b00;
			14'b00110000011100: M1r = 2'b00;
			14'b01110000011100: M1r = 2'b00;
			14'b10110000011100: M1r = 2'b00;
			14'b11110000011100: M1r = 2'b00;
			14'b00000100011100: M1r = 2'b00;
			14'b01000100011100: M1r = 2'b00;
			14'b10000100011100: M1r = 2'b00;
			14'b11000100011100: M1r = 2'b00;
			14'b00010100011100: M1r = 2'b00;
			14'b01010100011100: M1r = 2'b00;
			14'b10010100011100: M1r = 2'b00;
			14'b11010100011100: M1r = 2'b00;
			14'b00100100011100: M1r = 2'b00;
			14'b01100100011100: M1r = 2'b00;
			14'b10100100011100: M1r = 2'b00;
			14'b11100100011100: M1r = 2'b00;
			14'b00110100011100: M1r = 2'b00;
			14'b01110100011100: M1r = 2'b00;
			14'b10110100011100: M1r = 2'b00;
			14'b11110100011100: M1r = 2'b00;
			14'b00001000011100: M1r = 2'b00;
			14'b01001000011100: M1r = 2'b00;
			14'b10001000011100: M1r = 2'b00;
			14'b11001000011100: M1r = 2'b00;
			14'b00011000011100: M1r = 2'b00;
			14'b01011000011100: M1r = 2'b00;
			14'b10011000011100: M1r = 2'b00;
			14'b11011000011100: M1r = 2'b00;
			14'b00101000011100: M1r = 2'b00;
			14'b01101000011100: M1r = 2'b00;
			14'b10101000011100: M1r = 2'b00;
			14'b11101000011100: M1r = 2'b00;
			14'b00111000011100: M1r = 2'b00;
			14'b01111000011100: M1r = 2'b00;
			14'b10111000011100: M1r = 2'b00;
			14'b11111000011100: M1r = 2'b00;
			14'b00001100011100: M1r = 2'b00;
			14'b01001100011100: M1r = 2'b00;
			14'b10001100011100: M1r = 2'b00;
			14'b11001100011100: M1r = 2'b00;
			14'b00011100011100: M1r = 2'b00;
			14'b01011100011100: M1r = 2'b00;
			14'b10011100011100: M1r = 2'b00;
			14'b11011100011100: M1r = 2'b00;
			14'b00101100011100: M1r = 2'b00;
			14'b01101100011100: M1r = 2'b00;
			14'b10101100011100: M1r = 2'b00;
			14'b11101100011100: M1r = 2'b00;
			14'b00111100011100: M1r = 2'b00;
			14'b01111100011100: M1r = 2'b00;
			14'b10111100011100: M1r = 2'b00;
			14'b11111100011100: M1r = 2'b00;
			14'b00000001011100: M1r = 2'b00;
			14'b01000001011100: M1r = 2'b00;
			14'b10000001011100: M1r = 2'b00;
			14'b11000001011100: M1r = 2'b00;
			14'b00010001011100: M1r = 2'b00;
			14'b01010001011100: M1r = 2'b00;
			14'b10010001011100: M1r = 2'b00;
			14'b11010001011100: M1r = 2'b00;
			14'b00100001011100: M1r = 2'b00;
			14'b01100001011100: M1r = 2'b00;
			14'b10100001011100: M1r = 2'b00;
			14'b11100001011100: M1r = 2'b00;
			14'b00110001011100: M1r = 2'b00;
			14'b01110001011100: M1r = 2'b00;
			14'b10110001011100: M1r = 2'b00;
			14'b11110001011100: M1r = 2'b00;
			14'b00000101011100: M1r = 2'b00;
			14'b01000101011100: M1r = 2'b00;
			14'b10000101011100: M1r = 2'b00;
			14'b11000101011100: M1r = 2'b00;
			14'b00010101011100: M1r = 2'b00;
			14'b01010101011100: M1r = 2'b00;
			14'b10010101011100: M1r = 2'b00;
			14'b11010101011100: M1r = 2'b00;
			14'b00100101011100: M1r = 2'b00;
			14'b01100101011100: M1r = 2'b00;
			14'b10100101011100: M1r = 2'b00;
			14'b11100101011100: M1r = 2'b00;
			14'b00110101011100: M1r = 2'b00;
			14'b01110101011100: M1r = 2'b00;
			14'b10110101011100: M1r = 2'b00;
			14'b11110101011100: M1r = 2'b00;
			14'b00001001011100: M1r = 2'b00;
			14'b01001001011100: M1r = 2'b00;
			14'b10001001011100: M1r = 2'b00;
			14'b11001001011100: M1r = 2'b00;
			14'b00011001011100: M1r = 2'b00;
			14'b01011001011100: M1r = 2'b00;
			14'b10011001011100: M1r = 2'b00;
			14'b11011001011100: M1r = 2'b00;
			14'b00101001011100: M1r = 2'b00;
			14'b01101001011100: M1r = 2'b00;
			14'b10101001011100: M1r = 2'b00;
			14'b11101001011100: M1r = 2'b00;
			14'b00111001011100: M1r = 2'b00;
			14'b01111001011100: M1r = 2'b00;
			14'b10111001011100: M1r = 2'b00;
			14'b11111001011100: M1r = 2'b00;
			14'b00001101011100: M1r = 2'b00;
			14'b01001101011100: M1r = 2'b00;
			14'b10001101011100: M1r = 2'b00;
			14'b11001101011100: M1r = 2'b00;
			14'b00011101011100: M1r = 2'b00;
			14'b01011101011100: M1r = 2'b00;
			14'b10011101011100: M1r = 2'b00;
			14'b11011101011100: M1r = 2'b00;
			14'b00101101011100: M1r = 2'b00;
			14'b01101101011100: M1r = 2'b00;
			14'b10101101011100: M1r = 2'b00;
			14'b11101101011100: M1r = 2'b00;
			14'b00111101011100: M1r = 2'b00;
			14'b01111101011100: M1r = 2'b00;
			14'b10111101011100: M1r = 2'b00;
			14'b11111101011100: M1r = 2'b00;
			14'b00000010011100: M1r = 2'b00;
			14'b01000010011100: M1r = 2'b00;
			14'b10000010011100: M1r = 2'b00;
			14'b11000010011100: M1r = 2'b00;
			14'b00010010011100: M1r = 2'b00;
			14'b01010010011100: M1r = 2'b00;
			14'b10010010011100: M1r = 2'b00;
			14'b11010010011100: M1r = 2'b00;
			14'b00100010011100: M1r = 2'b00;
			14'b01100010011100: M1r = 2'b00;
			14'b10100010011100: M1r = 2'b00;
			14'b11100010011100: M1r = 2'b00;
			14'b00110010011100: M1r = 2'b00;
			14'b01110010011100: M1r = 2'b00;
			14'b10110010011100: M1r = 2'b00;
			14'b11110010011100: M1r = 2'b00;
			14'b00000110011100: M1r = 2'b00;
			14'b01000110011100: M1r = 2'b00;
			14'b10000110011100: M1r = 2'b00;
			14'b11000110011100: M1r = 2'b00;
			14'b00010110011100: M1r = 2'b00;
			14'b01010110011100: M1r = 2'b00;
			14'b10010110011100: M1r = 2'b00;
			14'b11010110011100: M1r = 2'b00;
			14'b00100110011100: M1r = 2'b00;
			14'b01100110011100: M1r = 2'b00;
			14'b10100110011100: M1r = 2'b00;
			14'b11100110011100: M1r = 2'b00;
			14'b00110110011100: M1r = 2'b00;
			14'b01110110011100: M1r = 2'b00;
			14'b10110110011100: M1r = 2'b00;
			14'b11110110011100: M1r = 2'b00;
			14'b00001010011100: M1r = 2'b00;
			14'b01001010011100: M1r = 2'b00;
			14'b10001010011100: M1r = 2'b00;
			14'b11001010011100: M1r = 2'b00;
			14'b00011010011100: M1r = 2'b00;
			14'b01011010011100: M1r = 2'b00;
			14'b10011010011100: M1r = 2'b00;
			14'b11011010011100: M1r = 2'b00;
			14'b00101010011100: M1r = 2'b00;
			14'b01101010011100: M1r = 2'b00;
			14'b10101010011100: M1r = 2'b00;
			14'b11101010011100: M1r = 2'b00;
			14'b00111010011100: M1r = 2'b00;
			14'b01111010011100: M1r = 2'b00;
			14'b10111010011100: M1r = 2'b00;
			14'b11111010011100: M1r = 2'b00;
			14'b00001110011100: M1r = 2'b00;
			14'b01001110011100: M1r = 2'b00;
			14'b10001110011100: M1r = 2'b00;
			14'b11001110011100: M1r = 2'b00;
			14'b00011110011100: M1r = 2'b00;
			14'b01011110011100: M1r = 2'b00;
			14'b10011110011100: M1r = 2'b00;
			14'b11011110011100: M1r = 2'b00;
			14'b00101110011100: M1r = 2'b00;
			14'b01101110011100: M1r = 2'b00;
			14'b10101110011100: M1r = 2'b00;
			14'b11101110011100: M1r = 2'b00;
			14'b00111110011100: M1r = 2'b00;
			14'b01111110011100: M1r = 2'b00;
			14'b10111110011100: M1r = 2'b00;
			14'b11111110011100: M1r = 2'b00;
			14'b00000011011100: M1r = 2'b00;
			14'b01000011011100: M1r = 2'b00;
			14'b10000011011100: M1r = 2'b00;
			14'b11000011011100: M1r = 2'b00;
			14'b00010011011100: M1r = 2'b00;
			14'b01010011011100: M1r = 2'b00;
			14'b10010011011100: M1r = 2'b00;
			14'b11010011011100: M1r = 2'b00;
			14'b00100011011100: M1r = 2'b00;
			14'b01100011011100: M1r = 2'b00;
			14'b10100011011100: M1r = 2'b00;
			14'b11100011011100: M1r = 2'b00;
			14'b00110011011100: M1r = 2'b00;
			14'b01110011011100: M1r = 2'b00;
			14'b10110011011100: M1r = 2'b00;
			14'b11110011011100: M1r = 2'b00;
			14'b00000111011100: M1r = 2'b00;
			14'b01000111011100: M1r = 2'b00;
			14'b10000111011100: M1r = 2'b00;
			14'b11000111011100: M1r = 2'b00;
			14'b00010111011100: M1r = 2'b00;
			14'b01010111011100: M1r = 2'b00;
			14'b10010111011100: M1r = 2'b00;
			14'b11010111011100: M1r = 2'b00;
			14'b00100111011100: M1r = 2'b00;
			14'b01100111011100: M1r = 2'b00;
			14'b10100111011100: M1r = 2'b00;
			14'b11100111011100: M1r = 2'b00;
			14'b00110111011100: M1r = 2'b00;
			14'b01110111011100: M1r = 2'b00;
			14'b10110111011100: M1r = 2'b00;
			14'b11110111011100: M1r = 2'b00;
			14'b00001011011100: M1r = 2'b00;
			14'b01001011011100: M1r = 2'b00;
			14'b10001011011100: M1r = 2'b00;
			14'b11001011011100: M1r = 2'b00;
			14'b00011011011100: M1r = 2'b00;
			14'b01011011011100: M1r = 2'b00;
			14'b10011011011100: M1r = 2'b00;
			14'b11011011011100: M1r = 2'b00;
			14'b00101011011100: M1r = 2'b00;
			14'b01101011011100: M1r = 2'b00;
			14'b10101011011100: M1r = 2'b00;
			14'b11101011011100: M1r = 2'b00;
			14'b00111011011100: M1r = 2'b00;
			14'b01111011011100: M1r = 2'b00;
			14'b10111011011100: M1r = 2'b00;
			14'b11111011011100: M1r = 2'b00;
			14'b00001111011100: M1r = 2'b00;
			14'b01001111011100: M1r = 2'b00;
			14'b10001111011100: M1r = 2'b00;
			14'b11001111011100: M1r = 2'b00;
			14'b00011111011100: M1r = 2'b00;
			14'b01011111011100: M1r = 2'b00;
			14'b10011111011100: M1r = 2'b00;
			14'b11011111011100: M1r = 2'b00;
			14'b00101111011100: M1r = 2'b00;
			14'b01101111011100: M1r = 2'b00;
			14'b10101111011100: M1r = 2'b00;
			14'b11101111011100: M1r = 2'b00;
			14'b00111111011100: M1r = 2'b00;
			14'b01111111011100: M1r = 2'b00;
			14'b10111111011100: M1r = 2'b00;
			14'b11111111011100: M1r = 2'b00;
			14'b00000000101100: M1r = 2'b00;
			14'b01000000101100: M1r = 2'b00;
			14'b10000000101100: M1r = 2'b00;
			14'b11000000101100: M1r = 2'b00;
			14'b00010000101100: M1r = 2'b00;
			14'b01010000101100: M1r = 2'b00;
			14'b10010000101100: M1r = 2'b00;
			14'b11010000101100: M1r = 2'b00;
			14'b00100000101100: M1r = 2'b00;
			14'b01100000101100: M1r = 2'b00;
			14'b10100000101100: M1r = 2'b00;
			14'b11100000101100: M1r = 2'b00;
			14'b00110000101100: M1r = 2'b00;
			14'b01110000101100: M1r = 2'b00;
			14'b10110000101100: M1r = 2'b00;
			14'b11110000101100: M1r = 2'b00;
			14'b00000100101100: M1r = 2'b00;
			14'b01000100101100: M1r = 2'b00;
			14'b10000100101100: M1r = 2'b00;
			14'b11000100101100: M1r = 2'b00;
			14'b00010100101100: M1r = 2'b00;
			14'b01010100101100: M1r = 2'b00;
			14'b10010100101100: M1r = 2'b00;
			14'b11010100101100: M1r = 2'b00;
			14'b00100100101100: M1r = 2'b00;
			14'b01100100101100: M1r = 2'b00;
			14'b10100100101100: M1r = 2'b00;
			14'b11100100101100: M1r = 2'b00;
			14'b00110100101100: M1r = 2'b00;
			14'b01110100101100: M1r = 2'b00;
			14'b10110100101100: M1r = 2'b00;
			14'b11110100101100: M1r = 2'b00;
			14'b00001000101100: M1r = 2'b00;
			14'b01001000101100: M1r = 2'b00;
			14'b10001000101100: M1r = 2'b00;
			14'b11001000101100: M1r = 2'b00;
			14'b00011000101100: M1r = 2'b00;
			14'b01011000101100: M1r = 2'b00;
			14'b10011000101100: M1r = 2'b00;
			14'b11011000101100: M1r = 2'b00;
			14'b00101000101100: M1r = 2'b00;
			14'b01101000101100: M1r = 2'b00;
			14'b10101000101100: M1r = 2'b00;
			14'b11101000101100: M1r = 2'b00;
			14'b00111000101100: M1r = 2'b00;
			14'b01111000101100: M1r = 2'b00;
			14'b10111000101100: M1r = 2'b00;
			14'b11111000101100: M1r = 2'b00;
			14'b00001100101100: M1r = 2'b00;
			14'b01001100101100: M1r = 2'b00;
			14'b10001100101100: M1r = 2'b00;
			14'b11001100101100: M1r = 2'b00;
			14'b00011100101100: M1r = 2'b00;
			14'b01011100101100: M1r = 2'b00;
			14'b10011100101100: M1r = 2'b00;
			14'b11011100101100: M1r = 2'b00;
			14'b00101100101100: M1r = 2'b00;
			14'b01101100101100: M1r = 2'b00;
			14'b10101100101100: M1r = 2'b00;
			14'b11101100101100: M1r = 2'b00;
			14'b00111100101100: M1r = 2'b00;
			14'b01111100101100: M1r = 2'b00;
			14'b10111100101100: M1r = 2'b00;
			14'b11111100101100: M1r = 2'b00;
			14'b00000001101100: M1r = 2'b00;
			14'b01000001101100: M1r = 2'b00;
			14'b10000001101100: M1r = 2'b00;
			14'b11000001101100: M1r = 2'b00;
			14'b00010001101100: M1r = 2'b00;
			14'b01010001101100: M1r = 2'b00;
			14'b10010001101100: M1r = 2'b00;
			14'b11010001101100: M1r = 2'b00;
			14'b00100001101100: M1r = 2'b00;
			14'b01100001101100: M1r = 2'b00;
			14'b10100001101100: M1r = 2'b00;
			14'b11100001101100: M1r = 2'b00;
			14'b00110001101100: M1r = 2'b00;
			14'b01110001101100: M1r = 2'b00;
			14'b10110001101100: M1r = 2'b00;
			14'b11110001101100: M1r = 2'b00;
			14'b00000101101100: M1r = 2'b00;
			14'b01000101101100: M1r = 2'b00;
			14'b10000101101100: M1r = 2'b00;
			14'b11000101101100: M1r = 2'b00;
			14'b00010101101100: M1r = 2'b00;
			14'b01010101101100: M1r = 2'b00;
			14'b10010101101100: M1r = 2'b00;
			14'b11010101101100: M1r = 2'b00;
			14'b00100101101100: M1r = 2'b00;
			14'b01100101101100: M1r = 2'b00;
			14'b10100101101100: M1r = 2'b00;
			14'b11100101101100: M1r = 2'b00;
			14'b00110101101100: M1r = 2'b00;
			14'b01110101101100: M1r = 2'b00;
			14'b10110101101100: M1r = 2'b00;
			14'b11110101101100: M1r = 2'b00;
			14'b00001001101100: M1r = 2'b00;
			14'b01001001101100: M1r = 2'b00;
			14'b10001001101100: M1r = 2'b00;
			14'b11001001101100: M1r = 2'b00;
			14'b00011001101100: M1r = 2'b00;
			14'b01011001101100: M1r = 2'b00;
			14'b10011001101100: M1r = 2'b00;
			14'b11011001101100: M1r = 2'b00;
			14'b00101001101100: M1r = 2'b00;
			14'b01101001101100: M1r = 2'b00;
			14'b10101001101100: M1r = 2'b00;
			14'b11101001101100: M1r = 2'b00;
			14'b00111001101100: M1r = 2'b00;
			14'b01111001101100: M1r = 2'b00;
			14'b10111001101100: M1r = 2'b00;
			14'b11111001101100: M1r = 2'b00;
			14'b00001101101100: M1r = 2'b00;
			14'b01001101101100: M1r = 2'b00;
			14'b10001101101100: M1r = 2'b00;
			14'b11001101101100: M1r = 2'b00;
			14'b00011101101100: M1r = 2'b00;
			14'b01011101101100: M1r = 2'b00;
			14'b10011101101100: M1r = 2'b00;
			14'b11011101101100: M1r = 2'b00;
			14'b00101101101100: M1r = 2'b00;
			14'b01101101101100: M1r = 2'b00;
			14'b10101101101100: M1r = 2'b00;
			14'b11101101101100: M1r = 2'b00;
			14'b00111101101100: M1r = 2'b00;
			14'b01111101101100: M1r = 2'b00;
			14'b10111101101100: M1r = 2'b00;
			14'b11111101101100: M1r = 2'b00;
			14'b00000010101100: M1r = 2'b00;
			14'b01000010101100: M1r = 2'b00;
			14'b10000010101100: M1r = 2'b00;
			14'b11000010101100: M1r = 2'b00;
			14'b00010010101100: M1r = 2'b00;
			14'b01010010101100: M1r = 2'b00;
			14'b10010010101100: M1r = 2'b00;
			14'b11010010101100: M1r = 2'b00;
			14'b00100010101100: M1r = 2'b00;
			14'b01100010101100: M1r = 2'b00;
			14'b10100010101100: M1r = 2'b00;
			14'b11100010101100: M1r = 2'b00;
			14'b00110010101100: M1r = 2'b00;
			14'b01110010101100: M1r = 2'b00;
			14'b10110010101100: M1r = 2'b00;
			14'b11110010101100: M1r = 2'b00;
			14'b00000110101100: M1r = 2'b00;
			14'b01000110101100: M1r = 2'b00;
			14'b10000110101100: M1r = 2'b00;
			14'b11000110101100: M1r = 2'b00;
			14'b00010110101100: M1r = 2'b00;
			14'b01010110101100: M1r = 2'b00;
			14'b10010110101100: M1r = 2'b00;
			14'b11010110101100: M1r = 2'b00;
			14'b00100110101100: M1r = 2'b00;
			14'b01100110101100: M1r = 2'b00;
			14'b10100110101100: M1r = 2'b00;
			14'b11100110101100: M1r = 2'b00;
			14'b00110110101100: M1r = 2'b00;
			14'b01110110101100: M1r = 2'b00;
			14'b10110110101100: M1r = 2'b00;
			14'b11110110101100: M1r = 2'b00;
			14'b00001010101100: M1r = 2'b00;
			14'b01001010101100: M1r = 2'b00;
			14'b10001010101100: M1r = 2'b00;
			14'b11001010101100: M1r = 2'b00;
			14'b00011010101100: M1r = 2'b00;
			14'b01011010101100: M1r = 2'b00;
			14'b10011010101100: M1r = 2'b00;
			14'b11011010101100: M1r = 2'b00;
			14'b00101010101100: M1r = 2'b00;
			14'b01101010101100: M1r = 2'b00;
			14'b10101010101100: M1r = 2'b00;
			14'b11101010101100: M1r = 2'b00;
			14'b00111010101100: M1r = 2'b00;
			14'b01111010101100: M1r = 2'b00;
			14'b10111010101100: M1r = 2'b00;
			14'b11111010101100: M1r = 2'b00;
			14'b00001110101100: M1r = 2'b00;
			14'b01001110101100: M1r = 2'b00;
			14'b10001110101100: M1r = 2'b00;
			14'b11001110101100: M1r = 2'b00;
			14'b00011110101100: M1r = 2'b00;
			14'b01011110101100: M1r = 2'b00;
			14'b10011110101100: M1r = 2'b00;
			14'b11011110101100: M1r = 2'b00;
			14'b00101110101100: M1r = 2'b00;
			14'b01101110101100: M1r = 2'b00;
			14'b10101110101100: M1r = 2'b00;
			14'b11101110101100: M1r = 2'b00;
			14'b00111110101100: M1r = 2'b00;
			14'b01111110101100: M1r = 2'b00;
			14'b10111110101100: M1r = 2'b00;
			14'b11111110101100: M1r = 2'b00;
			14'b00000011101100: M1r = 2'b00;
			14'b01000011101100: M1r = 2'b00;
			14'b10000011101100: M1r = 2'b00;
			14'b11000011101100: M1r = 2'b00;
			14'b00010011101100: M1r = 2'b00;
			14'b01010011101100: M1r = 2'b00;
			14'b10010011101100: M1r = 2'b00;
			14'b11010011101100: M1r = 2'b00;
			14'b00100011101100: M1r = 2'b00;
			14'b01100011101100: M1r = 2'b00;
			14'b10100011101100: M1r = 2'b00;
			14'b11100011101100: M1r = 2'b00;
			14'b00110011101100: M1r = 2'b00;
			14'b01110011101100: M1r = 2'b00;
			14'b10110011101100: M1r = 2'b00;
			14'b11110011101100: M1r = 2'b00;
			14'b00000111101100: M1r = 2'b00;
			14'b01000111101100: M1r = 2'b00;
			14'b10000111101100: M1r = 2'b00;
			14'b11000111101100: M1r = 2'b00;
			14'b00010111101100: M1r = 2'b00;
			14'b01010111101100: M1r = 2'b00;
			14'b10010111101100: M1r = 2'b00;
			14'b11010111101100: M1r = 2'b00;
			14'b00100111101100: M1r = 2'b00;
			14'b01100111101100: M1r = 2'b00;
			14'b10100111101100: M1r = 2'b00;
			14'b11100111101100: M1r = 2'b00;
			14'b00110111101100: M1r = 2'b00;
			14'b01110111101100: M1r = 2'b00;
			14'b10110111101100: M1r = 2'b00;
			14'b11110111101100: M1r = 2'b00;
			14'b00001011101100: M1r = 2'b00;
			14'b01001011101100: M1r = 2'b00;
			14'b10001011101100: M1r = 2'b00;
			14'b11001011101100: M1r = 2'b00;
			14'b00011011101100: M1r = 2'b00;
			14'b01011011101100: M1r = 2'b00;
			14'b10011011101100: M1r = 2'b00;
			14'b11011011101100: M1r = 2'b00;
			14'b00101011101100: M1r = 2'b00;
			14'b01101011101100: M1r = 2'b00;
			14'b10101011101100: M1r = 2'b00;
			14'b11101011101100: M1r = 2'b00;
			14'b00111011101100: M1r = 2'b00;
			14'b01111011101100: M1r = 2'b00;
			14'b10111011101100: M1r = 2'b00;
			14'b11111011101100: M1r = 2'b00;
			14'b00001111101100: M1r = 2'b00;
			14'b01001111101100: M1r = 2'b00;
			14'b10001111101100: M1r = 2'b00;
			14'b11001111101100: M1r = 2'b00;
			14'b00011111101100: M1r = 2'b00;
			14'b01011111101100: M1r = 2'b00;
			14'b10011111101100: M1r = 2'b00;
			14'b11011111101100: M1r = 2'b00;
			14'b00101111101100: M1r = 2'b00;
			14'b01101111101100: M1r = 2'b00;
			14'b10101111101100: M1r = 2'b00;
			14'b11101111101100: M1r = 2'b00;
			14'b00111111101100: M1r = 2'b00;
			14'b01111111101100: M1r = 2'b00;
			14'b10111111101100: M1r = 2'b00;
			14'b11111111101100: M1r = 2'b00;
			14'b00000000111100: M1r = 2'b00;
			14'b01000000111100: M1r = 2'b00;
			14'b10000000111100: M1r = 2'b00;
			14'b11000000111100: M1r = 2'b00;
			14'b00010000111100: M1r = 2'b00;
			14'b01010000111100: M1r = 2'b00;
			14'b10010000111100: M1r = 2'b00;
			14'b11010000111100: M1r = 2'b00;
			14'b00100000111100: M1r = 2'b00;
			14'b01100000111100: M1r = 2'b00;
			14'b10100000111100: M1r = 2'b00;
			14'b11100000111100: M1r = 2'b00;
			14'b00110000111100: M1r = 2'b00;
			14'b01110000111100: M1r = 2'b00;
			14'b10110000111100: M1r = 2'b00;
			14'b11110000111100: M1r = 2'b00;
			14'b00000100111100: M1r = 2'b00;
			14'b01000100111100: M1r = 2'b00;
			14'b10000100111100: M1r = 2'b00;
			14'b11000100111100: M1r = 2'b00;
			14'b00010100111100: M1r = 2'b00;
			14'b01010100111100: M1r = 2'b00;
			14'b10010100111100: M1r = 2'b00;
			14'b11010100111100: M1r = 2'b00;
			14'b00100100111100: M1r = 2'b00;
			14'b01100100111100: M1r = 2'b00;
			14'b10100100111100: M1r = 2'b00;
			14'b11100100111100: M1r = 2'b00;
			14'b00110100111100: M1r = 2'b00;
			14'b01110100111100: M1r = 2'b00;
			14'b10110100111100: M1r = 2'b00;
			14'b11110100111100: M1r = 2'b00;
			14'b00001000111100: M1r = 2'b00;
			14'b01001000111100: M1r = 2'b00;
			14'b10001000111100: M1r = 2'b00;
			14'b11001000111100: M1r = 2'b00;
			14'b00011000111100: M1r = 2'b00;
			14'b01011000111100: M1r = 2'b00;
			14'b10011000111100: M1r = 2'b00;
			14'b11011000111100: M1r = 2'b00;
			14'b00101000111100: M1r = 2'b00;
			14'b01101000111100: M1r = 2'b00;
			14'b10101000111100: M1r = 2'b00;
			14'b11101000111100: M1r = 2'b00;
			14'b00111000111100: M1r = 2'b00;
			14'b01111000111100: M1r = 2'b00;
			14'b10111000111100: M1r = 2'b00;
			14'b11111000111100: M1r = 2'b00;
			14'b00001100111100: M1r = 2'b00;
			14'b01001100111100: M1r = 2'b01;
			14'b10001100111100: M1r = 2'b01;
			14'b11001100111100: M1r = 2'b01;
			14'b00011100111100: M1r = 2'b00;
			14'b01011100111100: M1r = 2'b00;
			14'b10011100111100: M1r = 2'b00;
			14'b11011100111100: M1r = 2'b00;
			14'b00101100111100: M1r = 2'b00;
			14'b01101100111100: M1r = 2'b00;
			14'b10101100111100: M1r = 2'b00;
			14'b11101100111100: M1r = 2'b00;
			14'b00111100111100: M1r = 2'b00;
			14'b01111100111100: M1r = 2'b00;
			14'b10111100111100: M1r = 2'b00;
			14'b11111100111100: M1r = 2'b00;
			14'b00000001111100: M1r = 2'b00;
			14'b01000001111100: M1r = 2'b00;
			14'b10000001111100: M1r = 2'b00;
			14'b11000001111100: M1r = 2'b00;
			14'b00010001111100: M1r = 2'b00;
			14'b01010001111100: M1r = 2'b00;
			14'b10010001111100: M1r = 2'b00;
			14'b11010001111100: M1r = 2'b00;
			14'b00100001111100: M1r = 2'b00;
			14'b01100001111100: M1r = 2'b00;
			14'b10100001111100: M1r = 2'b00;
			14'b11100001111100: M1r = 2'b00;
			14'b00110001111100: M1r = 2'b00;
			14'b01110001111100: M1r = 2'b00;
			14'b10110001111100: M1r = 2'b00;
			14'b11110001111100: M1r = 2'b00;
			14'b00000101111100: M1r = 2'b00;
			14'b01000101111100: M1r = 2'b00;
			14'b10000101111100: M1r = 2'b00;
			14'b11000101111100: M1r = 2'b00;
			14'b00010101111100: M1r = 2'b00;
			14'b01010101111100: M1r = 2'b00;
			14'b10010101111100: M1r = 2'b00;
			14'b11010101111100: M1r = 2'b00;
			14'b00100101111100: M1r = 2'b00;
			14'b01100101111100: M1r = 2'b00;
			14'b10100101111100: M1r = 2'b00;
			14'b11100101111100: M1r = 2'b00;
			14'b00110101111100: M1r = 2'b00;
			14'b01110101111100: M1r = 2'b00;
			14'b10110101111100: M1r = 2'b00;
			14'b11110101111100: M1r = 2'b00;
			14'b00001001111100: M1r = 2'b00;
			14'b01001001111100: M1r = 2'b00;
			14'b10001001111100: M1r = 2'b00;
			14'b11001001111100: M1r = 2'b00;
			14'b00011001111100: M1r = 2'b00;
			14'b01011001111100: M1r = 2'b00;
			14'b10011001111100: M1r = 2'b00;
			14'b11011001111100: M1r = 2'b00;
			14'b00101001111100: M1r = 2'b00;
			14'b01101001111100: M1r = 2'b00;
			14'b10101001111100: M1r = 2'b00;
			14'b11101001111100: M1r = 2'b00;
			14'b00111001111100: M1r = 2'b00;
			14'b01111001111100: M1r = 2'b00;
			14'b10111001111100: M1r = 2'b00;
			14'b11111001111100: M1r = 2'b00;
			14'b00001101111100: M1r = 2'b00;
			14'b01001101111100: M1r = 2'b00;
			14'b10001101111100: M1r = 2'b00;
			14'b11001101111100: M1r = 2'b01;
			14'b00011101111100: M1r = 2'b00;
			14'b01011101111100: M1r = 2'b00;
			14'b10011101111100: M1r = 2'b00;
			14'b11011101111100: M1r = 2'b00;
			14'b00101101111100: M1r = 2'b00;
			14'b01101101111100: M1r = 2'b00;
			14'b10101101111100: M1r = 2'b00;
			14'b11101101111100: M1r = 2'b00;
			14'b00111101111100: M1r = 2'b00;
			14'b01111101111100: M1r = 2'b00;
			14'b10111101111100: M1r = 2'b00;
			14'b11111101111100: M1r = 2'b00;
			14'b00000010111100: M1r = 2'b00;
			14'b01000010111100: M1r = 2'b00;
			14'b10000010111100: M1r = 2'b00;
			14'b11000010111100: M1r = 2'b00;
			14'b00010010111100: M1r = 2'b00;
			14'b01010010111100: M1r = 2'b00;
			14'b10010010111100: M1r = 2'b00;
			14'b11010010111100: M1r = 2'b00;
			14'b00100010111100: M1r = 2'b00;
			14'b01100010111100: M1r = 2'b00;
			14'b10100010111100: M1r = 2'b00;
			14'b11100010111100: M1r = 2'b00;
			14'b00110010111100: M1r = 2'b00;
			14'b01110010111100: M1r = 2'b00;
			14'b10110010111100: M1r = 2'b00;
			14'b11110010111100: M1r = 2'b00;
			14'b00000110111100: M1r = 2'b00;
			14'b01000110111100: M1r = 2'b00;
			14'b10000110111100: M1r = 2'b00;
			14'b11000110111100: M1r = 2'b00;
			14'b00010110111100: M1r = 2'b00;
			14'b01010110111100: M1r = 2'b00;
			14'b10010110111100: M1r = 2'b00;
			14'b11010110111100: M1r = 2'b00;
			14'b00100110111100: M1r = 2'b00;
			14'b01100110111100: M1r = 2'b00;
			14'b10100110111100: M1r = 2'b00;
			14'b11100110111100: M1r = 2'b00;
			14'b00110110111100: M1r = 2'b00;
			14'b01110110111100: M1r = 2'b00;
			14'b10110110111100: M1r = 2'b00;
			14'b11110110111100: M1r = 2'b00;
			14'b00001010111100: M1r = 2'b00;
			14'b01001010111100: M1r = 2'b00;
			14'b10001010111100: M1r = 2'b00;
			14'b11001010111100: M1r = 2'b00;
			14'b00011010111100: M1r = 2'b00;
			14'b01011010111100: M1r = 2'b00;
			14'b10011010111100: M1r = 2'b00;
			14'b11011010111100: M1r = 2'b00;
			14'b00101010111100: M1r = 2'b00;
			14'b01101010111100: M1r = 2'b00;
			14'b10101010111100: M1r = 2'b00;
			14'b11101010111100: M1r = 2'b00;
			14'b00111010111100: M1r = 2'b00;
			14'b01111010111100: M1r = 2'b00;
			14'b10111010111100: M1r = 2'b00;
			14'b11111010111100: M1r = 2'b00;
			14'b00001110111100: M1r = 2'b00;
			14'b01001110111100: M1r = 2'b00;
			14'b10001110111100: M1r = 2'b00;
			14'b11001110111100: M1r = 2'b00;
			14'b00011110111100: M1r = 2'b00;
			14'b01011110111100: M1r = 2'b00;
			14'b10011110111100: M1r = 2'b00;
			14'b11011110111100: M1r = 2'b00;
			14'b00101110111100: M1r = 2'b00;
			14'b01101110111100: M1r = 2'b00;
			14'b10101110111100: M1r = 2'b00;
			14'b11101110111100: M1r = 2'b00;
			14'b00111110111100: M1r = 2'b00;
			14'b01111110111100: M1r = 2'b00;
			14'b10111110111100: M1r = 2'b00;
			14'b11111110111100: M1r = 2'b00;
			14'b00000011111100: M1r = 2'b00;
			14'b01000011111100: M1r = 2'b00;
			14'b10000011111100: M1r = 2'b00;
			14'b11000011111100: M1r = 2'b00;
			14'b00010011111100: M1r = 2'b00;
			14'b01010011111100: M1r = 2'b00;
			14'b10010011111100: M1r = 2'b00;
			14'b11010011111100: M1r = 2'b00;
			14'b00100011111100: M1r = 2'b00;
			14'b01100011111100: M1r = 2'b00;
			14'b10100011111100: M1r = 2'b00;
			14'b11100011111100: M1r = 2'b00;
			14'b00110011111100: M1r = 2'b00;
			14'b01110011111100: M1r = 2'b00;
			14'b10110011111100: M1r = 2'b00;
			14'b11110011111100: M1r = 2'b00;
			14'b00000111111100: M1r = 2'b00;
			14'b01000111111100: M1r = 2'b00;
			14'b10000111111100: M1r = 2'b00;
			14'b11000111111100: M1r = 2'b00;
			14'b00010111111100: M1r = 2'b00;
			14'b01010111111100: M1r = 2'b00;
			14'b10010111111100: M1r = 2'b00;
			14'b11010111111100: M1r = 2'b00;
			14'b00100111111100: M1r = 2'b00;
			14'b01100111111100: M1r = 2'b00;
			14'b10100111111100: M1r = 2'b00;
			14'b11100111111100: M1r = 2'b00;
			14'b00110111111100: M1r = 2'b00;
			14'b01110111111100: M1r = 2'b00;
			14'b10110111111100: M1r = 2'b00;
			14'b11110111111100: M1r = 2'b00;
			14'b00001011111100: M1r = 2'b00;
			14'b01001011111100: M1r = 2'b00;
			14'b10001011111100: M1r = 2'b00;
			14'b11001011111100: M1r = 2'b00;
			14'b00011011111100: M1r = 2'b00;
			14'b01011011111100: M1r = 2'b00;
			14'b10011011111100: M1r = 2'b00;
			14'b11011011111100: M1r = 2'b00;
			14'b00101011111100: M1r = 2'b00;
			14'b01101011111100: M1r = 2'b00;
			14'b10101011111100: M1r = 2'b00;
			14'b11101011111100: M1r = 2'b00;
			14'b00111011111100: M1r = 2'b00;
			14'b01111011111100: M1r = 2'b00;
			14'b10111011111100: M1r = 2'b00;
			14'b11111011111100: M1r = 2'b00;
			14'b00001111111100: M1r = 2'b00;
			14'b01001111111100: M1r = 2'b00;
			14'b10001111111100: M1r = 2'b00;
			14'b11001111111100: M1r = 2'b00;
			14'b00011111111100: M1r = 2'b00;
			14'b01011111111100: M1r = 2'b00;
			14'b10011111111100: M1r = 2'b00;
			14'b11011111111100: M1r = 2'b00;
			14'b00101111111100: M1r = 2'b00;
			14'b01101111111100: M1r = 2'b00;
			14'b10101111111100: M1r = 2'b00;
			14'b11101111111100: M1r = 2'b00;
			14'b00111111111100: M1r = 2'b00;
			14'b01111111111100: M1r = 2'b00;
			14'b10111111111100: M1r = 2'b00;
			14'b11111111111100: M1r = 2'b00;
			14'b00000000000001: M1r = 2'b00;
			14'b01000000000001: M1r = 2'b00;
			14'b10000000000001: M1r = 2'b00;
			14'b11000000000001: M1r = 2'b01;
			14'b00010000000001: M1r = 2'b00;
			14'b01010000000001: M1r = 2'b00;
			14'b10010000000001: M1r = 2'b00;
			14'b11010000000001: M1r = 2'b00;
			14'b00100000000001: M1r = 2'b00;
			14'b01100000000001: M1r = 2'b00;
			14'b10100000000001: M1r = 2'b00;
			14'b11100000000001: M1r = 2'b00;
			14'b00110000000001: M1r = 2'b00;
			14'b01110000000001: M1r = 2'b00;
			14'b10110000000001: M1r = 2'b00;
			14'b11110000000001: M1r = 2'b00;
			14'b00000100000001: M1r = 2'b01;
			14'b01000100000001: M1r = 2'b01;
			14'b10000100000001: M1r = 2'b01;
			14'b11000100000001: M1r = 2'b01;
			14'b00010100000001: M1r = 2'b00;
			14'b01010100000001: M1r = 2'b01;
			14'b10010100000001: M1r = 2'b01;
			14'b11010100000001: M1r = 2'b01;
			14'b00100100000001: M1r = 2'b00;
			14'b01100100000001: M1r = 2'b00;
			14'b10100100000001: M1r = 2'b00;
			14'b11100100000001: M1r = 2'b00;
			14'b00110100000001: M1r = 2'b00;
			14'b01110100000001: M1r = 2'b00;
			14'b10110100000001: M1r = 2'b00;
			14'b11110100000001: M1r = 2'b00;
			14'b00001000000001: M1r = 2'b10;
			14'b01001000000001: M1r = 2'b10;
			14'b10001000000001: M1r = 2'b10;
			14'b11001000000001: M1r = 2'b10;
			14'b00011000000001: M1r = 2'b01;
			14'b01011000000001: M1r = 2'b01;
			14'b10011000000001: M1r = 2'b01;
			14'b11011000000001: M1r = 2'b10;
			14'b00101000000001: M1r = 2'b01;
			14'b01101000000001: M1r = 2'b01;
			14'b10101000000001: M1r = 2'b01;
			14'b11101000000001: M1r = 2'b01;
			14'b00111000000001: M1r = 2'b00;
			14'b01111000000001: M1r = 2'b00;
			14'b10111000000001: M1r = 2'b00;
			14'b11111000000001: M1r = 2'b01;
			14'b00001100000001: M1r = 2'b10;
			14'b01001100000001: M1r = 2'b11;
			14'b10001100000001: M1r = 2'b11;
			14'b11001100000001: M1r = 2'b11;
			14'b00011100000001: M1r = 2'b10;
			14'b01011100000001: M1r = 2'b10;
			14'b10011100000001: M1r = 2'b10;
			14'b11011100000001: M1r = 2'b10;
			14'b00101100000001: M1r = 2'b01;
			14'b01101100000001: M1r = 2'b10;
			14'b10101100000001: M1r = 2'b10;
			14'b11101100000001: M1r = 2'b10;
			14'b00111100000001: M1r = 2'b01;
			14'b01111100000001: M1r = 2'b01;
			14'b10111100000001: M1r = 2'b01;
			14'b11111100000001: M1r = 2'b01;
			14'b00000001000001: M1r = 2'b00;
			14'b01000001000001: M1r = 2'b00;
			14'b10000001000001: M1r = 2'b00;
			14'b11000001000001: M1r = 2'b00;
			14'b00010001000001: M1r = 2'b00;
			14'b01010001000001: M1r = 2'b00;
			14'b10010001000001: M1r = 2'b00;
			14'b11010001000001: M1r = 2'b00;
			14'b00100001000001: M1r = 2'b00;
			14'b01100001000001: M1r = 2'b00;
			14'b10100001000001: M1r = 2'b00;
			14'b11100001000001: M1r = 2'b00;
			14'b00110001000001: M1r = 2'b00;
			14'b01110001000001: M1r = 2'b00;
			14'b10110001000001: M1r = 2'b00;
			14'b11110001000001: M1r = 2'b00;
			14'b00000101000001: M1r = 2'b01;
			14'b01000101000001: M1r = 2'b01;
			14'b10000101000001: M1r = 2'b01;
			14'b11000101000001: M1r = 2'b01;
			14'b00010101000001: M1r = 2'b00;
			14'b01010101000001: M1r = 2'b00;
			14'b10010101000001: M1r = 2'b00;
			14'b11010101000001: M1r = 2'b01;
			14'b00100101000001: M1r = 2'b00;
			14'b01100101000001: M1r = 2'b00;
			14'b10100101000001: M1r = 2'b00;
			14'b11100101000001: M1r = 2'b00;
			14'b00110101000001: M1r = 2'b00;
			14'b01110101000001: M1r = 2'b00;
			14'b10110101000001: M1r = 2'b00;
			14'b11110101000001: M1r = 2'b00;
			14'b00001001000001: M1r = 2'b01;
			14'b01001001000001: M1r = 2'b01;
			14'b10001001000001: M1r = 2'b10;
			14'b11001001000001: M1r = 2'b10;
			14'b00011001000001: M1r = 2'b01;
			14'b01011001000001: M1r = 2'b01;
			14'b10011001000001: M1r = 2'b01;
			14'b11011001000001: M1r = 2'b01;
			14'b00101001000001: M1r = 2'b00;
			14'b01101001000001: M1r = 2'b01;
			14'b10101001000001: M1r = 2'b01;
			14'b11101001000001: M1r = 2'b01;
			14'b00111001000001: M1r = 2'b00;
			14'b01111001000001: M1r = 2'b00;
			14'b10111001000001: M1r = 2'b00;
			14'b11111001000001: M1r = 2'b00;
			14'b00001101000001: M1r = 2'b10;
			14'b01001101000001: M1r = 2'b10;
			14'b10001101000001: M1r = 2'b10;
			14'b11001101000001: M1r = 2'b11;
			14'b00011101000001: M1r = 2'b10;
			14'b01011101000001: M1r = 2'b10;
			14'b10011101000001: M1r = 2'b10;
			14'b11011101000001: M1r = 2'b10;
			14'b00101101000001: M1r = 2'b01;
			14'b01101101000001: M1r = 2'b01;
			14'b10101101000001: M1r = 2'b01;
			14'b11101101000001: M1r = 2'b10;
			14'b00111101000001: M1r = 2'b01;
			14'b01111101000001: M1r = 2'b01;
			14'b10111101000001: M1r = 2'b01;
			14'b11111101000001: M1r = 2'b01;
			14'b00000010000001: M1r = 2'b00;
			14'b01000010000001: M1r = 2'b00;
			14'b10000010000001: M1r = 2'b00;
			14'b11000010000001: M1r = 2'b00;
			14'b00010010000001: M1r = 2'b00;
			14'b01010010000001: M1r = 2'b00;
			14'b10010010000001: M1r = 2'b00;
			14'b11010010000001: M1r = 2'b00;
			14'b00100010000001: M1r = 2'b00;
			14'b01100010000001: M1r = 2'b00;
			14'b10100010000001: M1r = 2'b00;
			14'b11100010000001: M1r = 2'b00;
			14'b00110010000001: M1r = 2'b00;
			14'b01110010000001: M1r = 2'b00;
			14'b10110010000001: M1r = 2'b00;
			14'b11110010000001: M1r = 2'b00;
			14'b00000110000001: M1r = 2'b00;
			14'b01000110000001: M1r = 2'b00;
			14'b10000110000001: M1r = 2'b01;
			14'b11000110000001: M1r = 2'b01;
			14'b00010110000001: M1r = 2'b00;
			14'b01010110000001: M1r = 2'b00;
			14'b10010110000001: M1r = 2'b00;
			14'b11010110000001: M1r = 2'b00;
			14'b00100110000001: M1r = 2'b00;
			14'b01100110000001: M1r = 2'b00;
			14'b10100110000001: M1r = 2'b00;
			14'b11100110000001: M1r = 2'b00;
			14'b00110110000001: M1r = 2'b00;
			14'b01110110000001: M1r = 2'b00;
			14'b10110110000001: M1r = 2'b00;
			14'b11110110000001: M1r = 2'b00;
			14'b00001010000001: M1r = 2'b01;
			14'b01001010000001: M1r = 2'b01;
			14'b10001010000001: M1r = 2'b01;
			14'b11001010000001: M1r = 2'b10;
			14'b00011010000001: M1r = 2'b01;
			14'b01011010000001: M1r = 2'b01;
			14'b10011010000001: M1r = 2'b01;
			14'b11011010000001: M1r = 2'b01;
			14'b00101010000001: M1r = 2'b00;
			14'b01101010000001: M1r = 2'b00;
			14'b10101010000001: M1r = 2'b00;
			14'b11101010000001: M1r = 2'b01;
			14'b00111010000001: M1r = 2'b00;
			14'b01111010000001: M1r = 2'b00;
			14'b10111010000001: M1r = 2'b00;
			14'b11111010000001: M1r = 2'b00;
			14'b00001110000001: M1r = 2'b10;
			14'b01001110000001: M1r = 2'b10;
			14'b10001110000001: M1r = 2'b10;
			14'b11001110000001: M1r = 2'b10;
			14'b00011110000001: M1r = 2'b01;
			14'b01011110000001: M1r = 2'b01;
			14'b10011110000001: M1r = 2'b10;
			14'b11011110000001: M1r = 2'b10;
			14'b00101110000001: M1r = 2'b01;
			14'b01101110000001: M1r = 2'b01;
			14'b10101110000001: M1r = 2'b01;
			14'b11101110000001: M1r = 2'b01;
			14'b00111110000001: M1r = 2'b00;
			14'b01111110000001: M1r = 2'b01;
			14'b10111110000001: M1r = 2'b01;
			14'b11111110000001: M1r = 2'b01;
			14'b00000011000001: M1r = 2'b00;
			14'b01000011000001: M1r = 2'b00;
			14'b10000011000001: M1r = 2'b00;
			14'b11000011000001: M1r = 2'b00;
			14'b00010011000001: M1r = 2'b00;
			14'b01010011000001: M1r = 2'b00;
			14'b10010011000001: M1r = 2'b00;
			14'b11010011000001: M1r = 2'b00;
			14'b00100011000001: M1r = 2'b00;
			14'b01100011000001: M1r = 2'b00;
			14'b10100011000001: M1r = 2'b00;
			14'b11100011000001: M1r = 2'b00;
			14'b00110011000001: M1r = 2'b00;
			14'b01110011000001: M1r = 2'b00;
			14'b10110011000001: M1r = 2'b00;
			14'b11110011000001: M1r = 2'b00;
			14'b00000111000001: M1r = 2'b00;
			14'b01000111000001: M1r = 2'b00;
			14'b10000111000001: M1r = 2'b00;
			14'b11000111000001: M1r = 2'b00;
			14'b00010111000001: M1r = 2'b00;
			14'b01010111000001: M1r = 2'b00;
			14'b10010111000001: M1r = 2'b00;
			14'b11010111000001: M1r = 2'b00;
			14'b00100111000001: M1r = 2'b00;
			14'b01100111000001: M1r = 2'b00;
			14'b10100111000001: M1r = 2'b00;
			14'b11100111000001: M1r = 2'b00;
			14'b00110111000001: M1r = 2'b00;
			14'b01110111000001: M1r = 2'b00;
			14'b10110111000001: M1r = 2'b00;
			14'b11110111000001: M1r = 2'b00;
			14'b00001011000001: M1r = 2'b01;
			14'b01001011000001: M1r = 2'b01;
			14'b10001011000001: M1r = 2'b01;
			14'b11001011000001: M1r = 2'b01;
			14'b00011011000001: M1r = 2'b00;
			14'b01011011000001: M1r = 2'b00;
			14'b10011011000001: M1r = 2'b01;
			14'b11011011000001: M1r = 2'b01;
			14'b00101011000001: M1r = 2'b00;
			14'b01101011000001: M1r = 2'b00;
			14'b10101011000001: M1r = 2'b00;
			14'b11101011000001: M1r = 2'b00;
			14'b00111011000001: M1r = 2'b00;
			14'b01111011000001: M1r = 2'b00;
			14'b10111011000001: M1r = 2'b00;
			14'b11111011000001: M1r = 2'b00;
			14'b00001111000001: M1r = 2'b10;
			14'b01001111000001: M1r = 2'b10;
			14'b10001111000001: M1r = 2'b10;
			14'b11001111000001: M1r = 2'b10;
			14'b00011111000001: M1r = 2'b01;
			14'b01011111000001: M1r = 2'b01;
			14'b10011111000001: M1r = 2'b01;
			14'b11011111000001: M1r = 2'b10;
			14'b00101111000001: M1r = 2'b01;
			14'b01101111000001: M1r = 2'b01;
			14'b10101111000001: M1r = 2'b01;
			14'b11101111000001: M1r = 2'b01;
			14'b00111111000001: M1r = 2'b00;
			14'b01111111000001: M1r = 2'b00;
			14'b10111111000001: M1r = 2'b00;
			14'b11111111000001: M1r = 2'b01;
			14'b00000000010001: M1r = 2'b01;
			14'b01000000010001: M1r = 2'b01;
			14'b10000000010001: M1r = 2'b01;
			14'b11000000010001: M1r = 2'b01;
			14'b00010000010001: M1r = 2'b00;
			14'b01010000010001: M1r = 2'b00;
			14'b10010000010001: M1r = 2'b00;
			14'b11010000010001: M1r = 2'b01;
			14'b00100000010001: M1r = 2'b00;
			14'b01100000010001: M1r = 2'b00;
			14'b10100000010001: M1r = 2'b00;
			14'b11100000010001: M1r = 2'b00;
			14'b00110000010001: M1r = 2'b00;
			14'b01110000010001: M1r = 2'b00;
			14'b10110000010001: M1r = 2'b00;
			14'b11110000010001: M1r = 2'b00;
			14'b00000100010001: M1r = 2'b01;
			14'b01000100010001: M1r = 2'b01;
			14'b10000100010001: M1r = 2'b10;
			14'b11000100010001: M1r = 2'b10;
			14'b00010100010001: M1r = 2'b01;
			14'b01010100010001: M1r = 2'b01;
			14'b10010100010001: M1r = 2'b01;
			14'b11010100010001: M1r = 2'b01;
			14'b00100100010001: M1r = 2'b00;
			14'b01100100010001: M1r = 2'b00;
			14'b10100100010001: M1r = 2'b01;
			14'b11100100010001: M1r = 2'b01;
			14'b00110100010001: M1r = 2'b00;
			14'b01110100010001: M1r = 2'b00;
			14'b10110100010001: M1r = 2'b00;
			14'b11110100010001: M1r = 2'b00;
			14'b00001000010001: M1r = 2'b10;
			14'b01001000010001: M1r = 2'b10;
			14'b10001000010001: M1r = 2'b10;
			14'b11001000010001: M1r = 2'b10;
			14'b00011000010001: M1r = 2'b10;
			14'b01011000010001: M1r = 2'b10;
			14'b10011000010001: M1r = 2'b10;
			14'b11011000010001: M1r = 2'b10;
			14'b00101000010001: M1r = 2'b01;
			14'b01101000010001: M1r = 2'b01;
			14'b10101000010001: M1r = 2'b01;
			14'b11101000010001: M1r = 2'b10;
			14'b00111000010001: M1r = 2'b01;
			14'b01111000010001: M1r = 2'b01;
			14'b10111000010001: M1r = 2'b01;
			14'b11111000010001: M1r = 2'b01;
			14'b00001100010001: M1r = 2'b11;
			14'b01001100010001: M1r = 2'b11;
			14'b10001100010001: M1r = 2'b11;
			14'b11001100010001: M1r = 2'b11;
			14'b00011100010001: M1r = 2'b10;
			14'b01011100010001: M1r = 2'b10;
			14'b10011100010001: M1r = 2'b11;
			14'b11011100010001: M1r = 2'b11;
			14'b00101100010001: M1r = 2'b10;
			14'b01101100010001: M1r = 2'b10;
			14'b10101100010001: M1r = 2'b10;
			14'b11101100010001: M1r = 2'b10;
			14'b00111100010001: M1r = 2'b01;
			14'b01111100010001: M1r = 2'b10;
			14'b10111100010001: M1r = 2'b10;
			14'b11111100010001: M1r = 2'b10;
			14'b00000001010001: M1r = 2'b00;
			14'b01000001010001: M1r = 2'b00;
			14'b10000001010001: M1r = 2'b01;
			14'b11000001010001: M1r = 2'b01;
			14'b00010001010001: M1r = 2'b00;
			14'b01010001010001: M1r = 2'b00;
			14'b10010001010001: M1r = 2'b00;
			14'b11010001010001: M1r = 2'b00;
			14'b00100001010001: M1r = 2'b00;
			14'b01100001010001: M1r = 2'b00;
			14'b10100001010001: M1r = 2'b00;
			14'b11100001010001: M1r = 2'b00;
			14'b00110001010001: M1r = 2'b00;
			14'b01110001010001: M1r = 2'b00;
			14'b10110001010001: M1r = 2'b00;
			14'b11110001010001: M1r = 2'b00;
			14'b00000101010001: M1r = 2'b01;
			14'b01000101010001: M1r = 2'b01;
			14'b10000101010001: M1r = 2'b01;
			14'b11000101010001: M1r = 2'b01;
			14'b00010101010001: M1r = 2'b01;
			14'b01010101010001: M1r = 2'b01;
			14'b10010101010001: M1r = 2'b01;
			14'b11010101010001: M1r = 2'b01;
			14'b00100101010001: M1r = 2'b00;
			14'b01100101010001: M1r = 2'b00;
			14'b10100101010001: M1r = 2'b00;
			14'b11100101010001: M1r = 2'b01;
			14'b00110101010001: M1r = 2'b00;
			14'b01110101010001: M1r = 2'b00;
			14'b10110101010001: M1r = 2'b00;
			14'b11110101010001: M1r = 2'b00;
			14'b00001001010001: M1r = 2'b10;
			14'b01001001010001: M1r = 2'b10;
			14'b10001001010001: M1r = 2'b10;
			14'b11001001010001: M1r = 2'b10;
			14'b00011001010001: M1r = 2'b01;
			14'b01011001010001: M1r = 2'b01;
			14'b10011001010001: M1r = 2'b10;
			14'b11011001010001: M1r = 2'b10;
			14'b00101001010001: M1r = 2'b01;
			14'b01101001010001: M1r = 2'b01;
			14'b10101001010001: M1r = 2'b01;
			14'b11101001010001: M1r = 2'b01;
			14'b00111001010001: M1r = 2'b00;
			14'b01111001010001: M1r = 2'b00;
			14'b10111001010001: M1r = 2'b01;
			14'b11111001010001: M1r = 2'b01;
			14'b00001101010001: M1r = 2'b11;
			14'b01001101010001: M1r = 2'b11;
			14'b10001101010001: M1r = 2'b11;
			14'b11001101010001: M1r = 2'b11;
			14'b00011101010001: M1r = 2'b10;
			14'b01011101010001: M1r = 2'b10;
			14'b10011101010001: M1r = 2'b10;
			14'b11011101010001: M1r = 2'b10;
			14'b00101101010001: M1r = 2'b10;
			14'b01101101010001: M1r = 2'b10;
			14'b10101101010001: M1r = 2'b10;
			14'b11101101010001: M1r = 2'b10;
			14'b00111101010001: M1r = 2'b01;
			14'b01111101010001: M1r = 2'b01;
			14'b10111101010001: M1r = 2'b01;
			14'b11111101010001: M1r = 2'b10;
			14'b00000010010001: M1r = 2'b00;
			14'b01000010010001: M1r = 2'b00;
			14'b10000010010001: M1r = 2'b00;
			14'b11000010010001: M1r = 2'b00;
			14'b00010010010001: M1r = 2'b00;
			14'b01010010010001: M1r = 2'b00;
			14'b10010010010001: M1r = 2'b00;
			14'b11010010010001: M1r = 2'b00;
			14'b00100010010001: M1r = 2'b00;
			14'b01100010010001: M1r = 2'b00;
			14'b10100010010001: M1r = 2'b00;
			14'b11100010010001: M1r = 2'b00;
			14'b00110010010001: M1r = 2'b00;
			14'b01110010010001: M1r = 2'b00;
			14'b10110010010001: M1r = 2'b00;
			14'b11110010010001: M1r = 2'b00;
			14'b00000110010001: M1r = 2'b01;
			14'b01000110010001: M1r = 2'b01;
			14'b10000110010001: M1r = 2'b01;
			14'b11000110010001: M1r = 2'b01;
			14'b00010110010001: M1r = 2'b00;
			14'b01010110010001: M1r = 2'b00;
			14'b10010110010001: M1r = 2'b01;
			14'b11010110010001: M1r = 2'b01;
			14'b00100110010001: M1r = 2'b00;
			14'b01100110010001: M1r = 2'b00;
			14'b10100110010001: M1r = 2'b00;
			14'b11100110010001: M1r = 2'b00;
			14'b00110110010001: M1r = 2'b00;
			14'b01110110010001: M1r = 2'b00;
			14'b10110110010001: M1r = 2'b00;
			14'b11110110010001: M1r = 2'b00;
			14'b00001010010001: M1r = 2'b01;
			14'b01001010010001: M1r = 2'b10;
			14'b10001010010001: M1r = 2'b10;
			14'b11001010010001: M1r = 2'b10;
			14'b00011010010001: M1r = 2'b01;
			14'b01011010010001: M1r = 2'b01;
			14'b10011010010001: M1r = 2'b01;
			14'b11011010010001: M1r = 2'b01;
			14'b00101010010001: M1r = 2'b01;
			14'b01101010010001: M1r = 2'b01;
			14'b10101010010001: M1r = 2'b01;
			14'b11101010010001: M1r = 2'b01;
			14'b00111010010001: M1r = 2'b00;
			14'b01111010010001: M1r = 2'b00;
			14'b10111010010001: M1r = 2'b00;
			14'b11111010010001: M1r = 2'b01;
			14'b00001110010001: M1r = 2'b10;
			14'b01001110010001: M1r = 2'b10;
			14'b10001110010001: M1r = 2'b11;
			14'b11001110010001: M1r = 2'b11;
			14'b00011110010001: M1r = 2'b10;
			14'b01011110010001: M1r = 2'b10;
			14'b10011110010001: M1r = 2'b10;
			14'b11011110010001: M1r = 2'b10;
			14'b00101110010001: M1r = 2'b01;
			14'b01101110010001: M1r = 2'b01;
			14'b10101110010001: M1r = 2'b10;
			14'b11101110010001: M1r = 2'b10;
			14'b00111110010001: M1r = 2'b01;
			14'b01111110010001: M1r = 2'b01;
			14'b10111110010001: M1r = 2'b01;
			14'b11111110010001: M1r = 2'b01;
			14'b00000011010001: M1r = 2'b00;
			14'b01000011010001: M1r = 2'b00;
			14'b10000011010001: M1r = 2'b00;
			14'b11000011010001: M1r = 2'b00;
			14'b00010011010001: M1r = 2'b00;
			14'b01010011010001: M1r = 2'b00;
			14'b10010011010001: M1r = 2'b00;
			14'b11010011010001: M1r = 2'b00;
			14'b00100011010001: M1r = 2'b00;
			14'b01100011010001: M1r = 2'b00;
			14'b10100011010001: M1r = 2'b00;
			14'b11100011010001: M1r = 2'b00;
			14'b00110011010001: M1r = 2'b00;
			14'b01110011010001: M1r = 2'b00;
			14'b10110011010001: M1r = 2'b00;
			14'b11110011010001: M1r = 2'b00;
			14'b00000111010001: M1r = 2'b00;
			14'b01000111010001: M1r = 2'b01;
			14'b10000111010001: M1r = 2'b01;
			14'b11000111010001: M1r = 2'b01;
			14'b00010111010001: M1r = 2'b00;
			14'b01010111010001: M1r = 2'b00;
			14'b10010111010001: M1r = 2'b00;
			14'b11010111010001: M1r = 2'b00;
			14'b00100111010001: M1r = 2'b00;
			14'b01100111010001: M1r = 2'b00;
			14'b10100111010001: M1r = 2'b00;
			14'b11100111010001: M1r = 2'b00;
			14'b00110111010001: M1r = 2'b00;
			14'b01110111010001: M1r = 2'b00;
			14'b10110111010001: M1r = 2'b00;
			14'b11110111010001: M1r = 2'b00;
			14'b00001011010001: M1r = 2'b01;
			14'b01001011010001: M1r = 2'b01;
			14'b10001011010001: M1r = 2'b10;
			14'b11001011010001: M1r = 2'b10;
			14'b00011011010001: M1r = 2'b01;
			14'b01011011010001: M1r = 2'b01;
			14'b10011011010001: M1r = 2'b01;
			14'b11011011010001: M1r = 2'b01;
			14'b00101011010001: M1r = 2'b00;
			14'b01101011010001: M1r = 2'b00;
			14'b10101011010001: M1r = 2'b01;
			14'b11101011010001: M1r = 2'b01;
			14'b00111011010001: M1r = 2'b00;
			14'b01111011010001: M1r = 2'b00;
			14'b10111011010001: M1r = 2'b00;
			14'b11111011010001: M1r = 2'b00;
			14'b00001111010001: M1r = 2'b10;
			14'b01001111010001: M1r = 2'b10;
			14'b10001111010001: M1r = 2'b10;
			14'b11001111010001: M1r = 2'b10;
			14'b00011111010001: M1r = 2'b01;
			14'b01011111010001: M1r = 2'b10;
			14'b10011111010001: M1r = 2'b10;
			14'b11011111010001: M1r = 2'b10;
			14'b00101111010001: M1r = 2'b01;
			14'b01101111010001: M1r = 2'b01;
			14'b10101111010001: M1r = 2'b01;
			14'b11101111010001: M1r = 2'b01;
			14'b00111111010001: M1r = 2'b01;
			14'b01111111010001: M1r = 2'b01;
			14'b10111111010001: M1r = 2'b01;
			14'b11111111010001: M1r = 2'b01;
			14'b00000000100001: M1r = 2'b01;
			14'b01000000100001: M1r = 2'b01;
			14'b10000000100001: M1r = 2'b01;
			14'b11000000100001: M1r = 2'b01;
			14'b00010000100001: M1r = 2'b00;
			14'b01010000100001: M1r = 2'b01;
			14'b10010000100001: M1r = 2'b01;
			14'b11010000100001: M1r = 2'b01;
			14'b00100000100001: M1r = 2'b00;
			14'b01100000100001: M1r = 2'b00;
			14'b10100000100001: M1r = 2'b00;
			14'b11100000100001: M1r = 2'b00;
			14'b00110000100001: M1r = 2'b00;
			14'b01110000100001: M1r = 2'b00;
			14'b10110000100001: M1r = 2'b00;
			14'b11110000100001: M1r = 2'b00;
			14'b00000100100001: M1r = 2'b10;
			14'b01000100100001: M1r = 2'b10;
			14'b10000100100001: M1r = 2'b10;
			14'b11000100100001: M1r = 2'b10;
			14'b00010100100001: M1r = 2'b01;
			14'b01010100100001: M1r = 2'b01;
			14'b10010100100001: M1r = 2'b10;
			14'b11010100100001: M1r = 2'b10;
			14'b00100100100001: M1r = 2'b01;
			14'b01100100100001: M1r = 2'b01;
			14'b10100100100001: M1r = 2'b01;
			14'b11100100100001: M1r = 2'b01;
			14'b00110100100001: M1r = 2'b00;
			14'b01110100100001: M1r = 2'b00;
			14'b10110100100001: M1r = 2'b01;
			14'b11110100100001: M1r = 2'b01;
			14'b00001000100001: M1r = 2'b10;
			14'b01001000100001: M1r = 2'b11;
			14'b10001000100001: M1r = 2'b11;
			14'b11001000100001: M1r = 2'b11;
			14'b00011000100001: M1r = 2'b10;
			14'b01011000100001: M1r = 2'b10;
			14'b10011000100001: M1r = 2'b10;
			14'b11011000100001: M1r = 2'b10;
			14'b00101000100001: M1r = 2'b10;
			14'b01101000100001: M1r = 2'b10;
			14'b10101000100001: M1r = 2'b10;
			14'b11101000100001: M1r = 2'b10;
			14'b00111000100001: M1r = 2'b01;
			14'b01111000100001: M1r = 2'b01;
			14'b10111000100001: M1r = 2'b01;
			14'b11111000100001: M1r = 2'b10;
			14'b00001100100001: M1r = 2'b11;
			14'b01001100100001: M1r = 2'b11;
			14'b10001100100001: M1r = 2'b11;
			14'b11001100100001: M1r = 2'b11;
			14'b00011100100001: M1r = 2'b11;
			14'b01011100100001: M1r = 2'b11;
			14'b10011100100001: M1r = 2'b11;
			14'b11011100100001: M1r = 2'b11;
			14'b00101100100001: M1r = 2'b10;
			14'b01101100100001: M1r = 2'b10;
			14'b10101100100001: M1r = 2'b11;
			14'b11101100100001: M1r = 2'b11;
			14'b00111100100001: M1r = 2'b10;
			14'b01111100100001: M1r = 2'b10;
			14'b10111100100001: M1r = 2'b10;
			14'b11111100100001: M1r = 2'b10;
			14'b00000001100001: M1r = 2'b01;
			14'b01000001100001: M1r = 2'b01;
			14'b10000001100001: M1r = 2'b01;
			14'b11000001100001: M1r = 2'b01;
			14'b00010001100001: M1r = 2'b00;
			14'b01010001100001: M1r = 2'b00;
			14'b10010001100001: M1r = 2'b01;
			14'b11010001100001: M1r = 2'b01;
			14'b00100001100001: M1r = 2'b00;
			14'b01100001100001: M1r = 2'b00;
			14'b10100001100001: M1r = 2'b00;
			14'b11100001100001: M1r = 2'b00;
			14'b00110001100001: M1r = 2'b00;
			14'b01110001100001: M1r = 2'b00;
			14'b10110001100001: M1r = 2'b00;
			14'b11110001100001: M1r = 2'b00;
			14'b00000101100001: M1r = 2'b01;
			14'b01000101100001: M1r = 2'b10;
			14'b10000101100001: M1r = 2'b10;
			14'b11000101100001: M1r = 2'b10;
			14'b00010101100001: M1r = 2'b01;
			14'b01010101100001: M1r = 2'b01;
			14'b10010101100001: M1r = 2'b01;
			14'b11010101100001: M1r = 2'b01;
			14'b00100101100001: M1r = 2'b00;
			14'b01100101100001: M1r = 2'b01;
			14'b10100101100001: M1r = 2'b01;
			14'b11100101100001: M1r = 2'b01;
			14'b00110101100001: M1r = 2'b00;
			14'b01110101100001: M1r = 2'b00;
			14'b10110101100001: M1r = 2'b00;
			14'b11110101100001: M1r = 2'b00;
			14'b00001001100001: M1r = 2'b10;
			14'b01001001100001: M1r = 2'b10;
			14'b10001001100001: M1r = 2'b10;
			14'b11001001100001: M1r = 2'b11;
			14'b00011001100001: M1r = 2'b10;
			14'b01011001100001: M1r = 2'b10;
			14'b10011001100001: M1r = 2'b10;
			14'b11011001100001: M1r = 2'b10;
			14'b00101001100001: M1r = 2'b01;
			14'b01101001100001: M1r = 2'b01;
			14'b10101001100001: M1r = 2'b10;
			14'b11101001100001: M1r = 2'b10;
			14'b00111001100001: M1r = 2'b01;
			14'b01111001100001: M1r = 2'b01;
			14'b10111001100001: M1r = 2'b01;
			14'b11111001100001: M1r = 2'b01;
			14'b00001101100001: M1r = 2'b11;
			14'b01001101100001: M1r = 2'b11;
			14'b10001101100001: M1r = 2'b11;
			14'b11001101100001: M1r = 2'b11;
			14'b00011101100001: M1r = 2'b10;
			14'b01011101100001: M1r = 2'b11;
			14'b10011101100001: M1r = 2'b11;
			14'b11011101100001: M1r = 2'b11;
			14'b00101101100001: M1r = 2'b10;
			14'b01101101100001: M1r = 2'b10;
			14'b10101101100001: M1r = 2'b10;
			14'b11101101100001: M1r = 2'b10;
			14'b00111101100001: M1r = 2'b10;
			14'b01111101100001: M1r = 2'b10;
			14'b10111101100001: M1r = 2'b10;
			14'b11111101100001: M1r = 2'b10;
			14'b00000010100001: M1r = 2'b00;
			14'b01000010100001: M1r = 2'b01;
			14'b10000010100001: M1r = 2'b01;
			14'b11000010100001: M1r = 2'b01;
			14'b00010010100001: M1r = 2'b00;
			14'b01010010100001: M1r = 2'b00;
			14'b10010010100001: M1r = 2'b00;
			14'b11010010100001: M1r = 2'b00;
			14'b00100010100001: M1r = 2'b00;
			14'b01100010100001: M1r = 2'b00;
			14'b10100010100001: M1r = 2'b00;
			14'b11100010100001: M1r = 2'b00;
			14'b00110010100001: M1r = 2'b00;
			14'b01110010100001: M1r = 2'b00;
			14'b10110010100001: M1r = 2'b00;
			14'b11110010100001: M1r = 2'b00;
			14'b00000110100001: M1r = 2'b01;
			14'b01000110100001: M1r = 2'b01;
			14'b10000110100001: M1r = 2'b01;
			14'b11000110100001: M1r = 2'b10;
			14'b00010110100001: M1r = 2'b01;
			14'b01010110100001: M1r = 2'b01;
			14'b10010110100001: M1r = 2'b01;
			14'b11010110100001: M1r = 2'b01;
			14'b00100110100001: M1r = 2'b00;
			14'b01100110100001: M1r = 2'b00;
			14'b10100110100001: M1r = 2'b01;
			14'b11100110100001: M1r = 2'b01;
			14'b00110110100001: M1r = 2'b00;
			14'b01110110100001: M1r = 2'b00;
			14'b10110110100001: M1r = 2'b00;
			14'b11110110100001: M1r = 2'b00;
			14'b00001010100001: M1r = 2'b10;
			14'b01001010100001: M1r = 2'b10;
			14'b10001010100001: M1r = 2'b10;
			14'b11001010100001: M1r = 2'b10;
			14'b00011010100001: M1r = 2'b01;
			14'b01011010100001: M1r = 2'b10;
			14'b10011010100001: M1r = 2'b10;
			14'b11011010100001: M1r = 2'b10;
			14'b00101010100001: M1r = 2'b01;
			14'b01101010100001: M1r = 2'b01;
			14'b10101010100001: M1r = 2'b01;
			14'b11101010100001: M1r = 2'b01;
			14'b00111010100001: M1r = 2'b00;
			14'b01111010100001: M1r = 2'b01;
			14'b10111010100001: M1r = 2'b01;
			14'b11111010100001: M1r = 2'b01;
			14'b00001110100001: M1r = 2'b11;
			14'b01001110100001: M1r = 2'b11;
			14'b10001110100001: M1r = 2'b11;
			14'b11001110100001: M1r = 2'b11;
			14'b00011110100001: M1r = 2'b10;
			14'b01011110100001: M1r = 2'b10;
			14'b10011110100001: M1r = 2'b10;
			14'b11011110100001: M1r = 2'b11;
			14'b00101110100001: M1r = 2'b10;
			14'b01101110100001: M1r = 2'b10;
			14'b10101110100001: M1r = 2'b10;
			14'b11101110100001: M1r = 2'b10;
			14'b00111110100001: M1r = 2'b01;
			14'b01111110100001: M1r = 2'b01;
			14'b10111110100001: M1r = 2'b10;
			14'b11111110100001: M1r = 2'b10;
			14'b00000011100001: M1r = 2'b00;
			14'b01000011100001: M1r = 2'b00;
			14'b10000011100001: M1r = 2'b00;
			14'b11000011100001: M1r = 2'b01;
			14'b00010011100001: M1r = 2'b00;
			14'b01010011100001: M1r = 2'b00;
			14'b10010011100001: M1r = 2'b00;
			14'b11010011100001: M1r = 2'b00;
			14'b00100011100001: M1r = 2'b00;
			14'b01100011100001: M1r = 2'b00;
			14'b10100011100001: M1r = 2'b00;
			14'b11100011100001: M1r = 2'b00;
			14'b00110011100001: M1r = 2'b00;
			14'b01110011100001: M1r = 2'b00;
			14'b10110011100001: M1r = 2'b00;
			14'b11110011100001: M1r = 2'b00;
			14'b00000111100001: M1r = 2'b01;
			14'b01000111100001: M1r = 2'b01;
			14'b10000111100001: M1r = 2'b01;
			14'b11000111100001: M1r = 2'b01;
			14'b00010111100001: M1r = 2'b00;
			14'b01010111100001: M1r = 2'b01;
			14'b10010111100001: M1r = 2'b01;
			14'b11010111100001: M1r = 2'b01;
			14'b00100111100001: M1r = 2'b00;
			14'b01100111100001: M1r = 2'b00;
			14'b10100111100001: M1r = 2'b00;
			14'b11100111100001: M1r = 2'b00;
			14'b00110111100001: M1r = 2'b00;
			14'b01110111100001: M1r = 2'b00;
			14'b10110111100001: M1r = 2'b00;
			14'b11110111100001: M1r = 2'b00;
			14'b00001011100001: M1r = 2'b10;
			14'b01001011100001: M1r = 2'b10;
			14'b10001011100001: M1r = 2'b10;
			14'b11001011100001: M1r = 2'b10;
			14'b00011011100001: M1r = 2'b01;
			14'b01011011100001: M1r = 2'b01;
			14'b10011011100001: M1r = 2'b01;
			14'b11011011100001: M1r = 2'b10;
			14'b00101011100001: M1r = 2'b01;
			14'b01101011100001: M1r = 2'b01;
			14'b10101011100001: M1r = 2'b01;
			14'b11101011100001: M1r = 2'b01;
			14'b00111011100001: M1r = 2'b00;
			14'b01111011100001: M1r = 2'b00;
			14'b10111011100001: M1r = 2'b01;
			14'b11111011100001: M1r = 2'b01;
			14'b00001111100001: M1r = 2'b10;
			14'b01001111100001: M1r = 2'b11;
			14'b10001111100001: M1r = 2'b11;
			14'b11001111100001: M1r = 2'b11;
			14'b00011111100001: M1r = 2'b10;
			14'b01011111100001: M1r = 2'b10;
			14'b10011111100001: M1r = 2'b10;
			14'b11011111100001: M1r = 2'b10;
			14'b00101111100001: M1r = 2'b01;
			14'b01101111100001: M1r = 2'b10;
			14'b10101111100001: M1r = 2'b10;
			14'b11101111100001: M1r = 2'b10;
			14'b00111111100001: M1r = 2'b01;
			14'b01111111100001: M1r = 2'b01;
			14'b10111111100001: M1r = 2'b01;
			14'b11111111100001: M1r = 2'b01;
			14'b00000000110001: M1r = 2'b01;
			14'b01000000110001: M1r = 2'b10;
			14'b10000000110001: M1r = 2'b10;
			14'b11000000110001: M1r = 2'b10;
			14'b00010000110001: M1r = 2'b01;
			14'b01010000110001: M1r = 2'b01;
			14'b10010000110001: M1r = 2'b01;
			14'b11010000110001: M1r = 2'b01;
			14'b00100000110001: M1r = 2'b00;
			14'b01100000110001: M1r = 2'b01;
			14'b10100000110001: M1r = 2'b01;
			14'b11100000110001: M1r = 2'b01;
			14'b00110000110001: M1r = 2'b00;
			14'b01110000110001: M1r = 2'b00;
			14'b10110000110001: M1r = 2'b00;
			14'b11110000110001: M1r = 2'b00;
			14'b00000100110001: M1r = 2'b10;
			14'b01000100110001: M1r = 2'b10;
			14'b10000100110001: M1r = 2'b10;
			14'b11000100110001: M1r = 2'b11;
			14'b00010100110001: M1r = 2'b10;
			14'b01010100110001: M1r = 2'b10;
			14'b10010100110001: M1r = 2'b10;
			14'b11010100110001: M1r = 2'b10;
			14'b00100100110001: M1r = 2'b01;
			14'b01100100110001: M1r = 2'b01;
			14'b10100100110001: M1r = 2'b10;
			14'b11100100110001: M1r = 2'b10;
			14'b00110100110001: M1r = 2'b01;
			14'b01110100110001: M1r = 2'b01;
			14'b10110100110001: M1r = 2'b01;
			14'b11110100110001: M1r = 2'b01;
			14'b00001000110001: M1r = 2'b11;
			14'b01001000110001: M1r = 2'b11;
			14'b10001000110001: M1r = 2'b11;
			14'b11001000110001: M1r = 2'b11;
			14'b00011000110001: M1r = 2'b10;
			14'b01011000110001: M1r = 2'b11;
			14'b10011000110001: M1r = 2'b11;
			14'b11011000110001: M1r = 2'b11;
			14'b00101000110001: M1r = 2'b10;
			14'b01101000110001: M1r = 2'b10;
			14'b10101000110001: M1r = 2'b10;
			14'b11101000110001: M1r = 2'b10;
			14'b00111000110001: M1r = 2'b01;
			14'b01111000110001: M1r = 2'b10;
			14'b10111000110001: M1r = 2'b10;
			14'b11111000110001: M1r = 2'b10;
			14'b00001100110001: M1r = 2'b11;
			14'b01001100110001: M1r = 2'b11;
			14'b10001100110001: M1r = 2'b11;
			14'b11001100110001: M1r = 2'b11;
			14'b00011100110001: M1r = 2'b11;
			14'b01011100110001: M1r = 2'b11;
			14'b10011100110001: M1r = 2'b11;
			14'b11011100110001: M1r = 2'b11;
			14'b00101100110001: M1r = 2'b11;
			14'b01101100110001: M1r = 2'b11;
			14'b10101100110001: M1r = 2'b11;
			14'b11101100110001: M1r = 2'b11;
			14'b00111100110001: M1r = 2'b10;
			14'b01111100110001: M1r = 2'b10;
			14'b10111100110001: M1r = 2'b11;
			14'b11111100110001: M1r = 2'b11;
			14'b00000001110001: M1r = 2'b01;
			14'b01000001110001: M1r = 2'b01;
			14'b10000001110001: M1r = 2'b01;
			14'b11000001110001: M1r = 2'b10;
			14'b00010001110001: M1r = 2'b01;
			14'b01010001110001: M1r = 2'b01;
			14'b10010001110001: M1r = 2'b01;
			14'b11010001110001: M1r = 2'b01;
			14'b00100001110001: M1r = 2'b00;
			14'b01100001110001: M1r = 2'b00;
			14'b10100001110001: M1r = 2'b00;
			14'b11100001110001: M1r = 2'b01;
			14'b00110001110001: M1r = 2'b00;
			14'b01110001110001: M1r = 2'b00;
			14'b10110001110001: M1r = 2'b00;
			14'b11110001110001: M1r = 2'b00;
			14'b00000101110001: M1r = 2'b10;
			14'b01000101110001: M1r = 2'b10;
			14'b10000101110001: M1r = 2'b10;
			14'b11000101110001: M1r = 2'b10;
			14'b00010101110001: M1r = 2'b01;
			14'b01010101110001: M1r = 2'b10;
			14'b10010101110001: M1r = 2'b10;
			14'b11010101110001: M1r = 2'b10;
			14'b00100101110001: M1r = 2'b01;
			14'b01100101110001: M1r = 2'b01;
			14'b10100101110001: M1r = 2'b01;
			14'b11100101110001: M1r = 2'b01;
			14'b00110101110001: M1r = 2'b00;
			14'b01110101110001: M1r = 2'b01;
			14'b10110101110001: M1r = 2'b01;
			14'b11110101110001: M1r = 2'b01;
			14'b00001001110001: M1r = 2'b11;
			14'b01001001110001: M1r = 2'b11;
			14'b10001001110001: M1r = 2'b11;
			14'b11001001110001: M1r = 2'b11;
			14'b00011001110001: M1r = 2'b10;
			14'b01011001110001: M1r = 2'b10;
			14'b10011001110001: M1r = 2'b10;
			14'b11011001110001: M1r = 2'b11;
			14'b00101001110001: M1r = 2'b10;
			14'b01101001110001: M1r = 2'b10;
			14'b10101001110001: M1r = 2'b10;
			14'b11101001110001: M1r = 2'b10;
			14'b00111001110001: M1r = 2'b01;
			14'b01111001110001: M1r = 2'b01;
			14'b10111001110001: M1r = 2'b10;
			14'b11111001110001: M1r = 2'b10;
			14'b00001101110001: M1r = 2'b11;
			14'b01001101110001: M1r = 2'b11;
			14'b10001101110001: M1r = 2'b11;
			14'b11001101110001: M1r = 2'b11;
			14'b00011101110001: M1r = 2'b11;
			14'b01011101110001: M1r = 2'b11;
			14'b10011101110001: M1r = 2'b11;
			14'b11011101110001: M1r = 2'b11;
			14'b00101101110001: M1r = 2'b10;
			14'b01101101110001: M1r = 2'b11;
			14'b10101101110001: M1r = 2'b11;
			14'b11101101110001: M1r = 2'b11;
			14'b00111101110001: M1r = 2'b10;
			14'b01111101110001: M1r = 2'b10;
			14'b10111101110001: M1r = 2'b10;
			14'b11111101110001: M1r = 2'b10;
			14'b00000010110001: M1r = 2'b01;
			14'b01000010110001: M1r = 2'b01;
			14'b10000010110001: M1r = 2'b01;
			14'b11000010110001: M1r = 2'b01;
			14'b00010010110001: M1r = 2'b00;
			14'b01010010110001: M1r = 2'b01;
			14'b10010010110001: M1r = 2'b01;
			14'b11010010110001: M1r = 2'b01;
			14'b00100010110001: M1r = 2'b00;
			14'b01100010110001: M1r = 2'b00;
			14'b10100010110001: M1r = 2'b00;
			14'b11100010110001: M1r = 2'b00;
			14'b00110010110001: M1r = 2'b00;
			14'b01110010110001: M1r = 2'b00;
			14'b10110010110001: M1r = 2'b00;
			14'b11110010110001: M1r = 2'b00;
			14'b00000110110001: M1r = 2'b10;
			14'b01000110110001: M1r = 2'b10;
			14'b10000110110001: M1r = 2'b10;
			14'b11000110110001: M1r = 2'b10;
			14'b00010110110001: M1r = 2'b01;
			14'b01010110110001: M1r = 2'b01;
			14'b10010110110001: M1r = 2'b01;
			14'b11010110110001: M1r = 2'b10;
			14'b00100110110001: M1r = 2'b01;
			14'b01100110110001: M1r = 2'b01;
			14'b10100110110001: M1r = 2'b01;
			14'b11100110110001: M1r = 2'b01;
			14'b00110110110001: M1r = 2'b00;
			14'b01110110110001: M1r = 2'b00;
			14'b10110110110001: M1r = 2'b00;
			14'b11110110110001: M1r = 2'b01;
			14'b00001010110001: M1r = 2'b10;
			14'b01001010110001: M1r = 2'b11;
			14'b10001010110001: M1r = 2'b11;
			14'b11001010110001: M1r = 2'b11;
			14'b00011010110001: M1r = 2'b10;
			14'b01011010110001: M1r = 2'b10;
			14'b10011010110001: M1r = 2'b10;
			14'b11011010110001: M1r = 2'b10;
			14'b00101010110001: M1r = 2'b01;
			14'b01101010110001: M1r = 2'b10;
			14'b10101010110001: M1r = 2'b10;
			14'b11101010110001: M1r = 2'b10;
			14'b00111010110001: M1r = 2'b01;
			14'b01111010110001: M1r = 2'b01;
			14'b10111010110001: M1r = 2'b01;
			14'b11111010110001: M1r = 2'b01;
			14'b00001110110001: M1r = 2'b11;
			14'b01001110110001: M1r = 2'b11;
			14'b10001110110001: M1r = 2'b11;
			14'b11001110110001: M1r = 2'b11;
			14'b00011110110001: M1r = 2'b11;
			14'b01011110110001: M1r = 2'b11;
			14'b10011110110001: M1r = 2'b11;
			14'b11011110110001: M1r = 2'b11;
			14'b00101110110001: M1r = 2'b10;
			14'b01101110110001: M1r = 2'b10;
			14'b10101110110001: M1r = 2'b10;
			14'b11101110110001: M1r = 2'b11;
			14'b00111110110001: M1r = 2'b10;
			14'b01111110110001: M1r = 2'b10;
			14'b10111110110001: M1r = 2'b10;
			14'b11111110110001: M1r = 2'b10;
			14'b00000011110001: M1r = 2'b01;
			14'b01000011110001: M1r = 2'b01;
			14'b10000011110001: M1r = 2'b01;
			14'b11000011110001: M1r = 2'b01;
			14'b00010011110001: M1r = 2'b00;
			14'b01010011110001: M1r = 2'b00;
			14'b10010011110001: M1r = 2'b00;
			14'b11010011110001: M1r = 2'b01;
			14'b00100011110001: M1r = 2'b00;
			14'b01100011110001: M1r = 2'b00;
			14'b10100011110001: M1r = 2'b00;
			14'b11100011110001: M1r = 2'b00;
			14'b00110011110001: M1r = 2'b00;
			14'b01110011110001: M1r = 2'b00;
			14'b10110011110001: M1r = 2'b00;
			14'b11110011110001: M1r = 2'b00;
			14'b00000111110001: M1r = 2'b01;
			14'b01000111110001: M1r = 2'b01;
			14'b10000111110001: M1r = 2'b10;
			14'b11000111110001: M1r = 2'b10;
			14'b00010111110001: M1r = 2'b01;
			14'b01010111110001: M1r = 2'b01;
			14'b10010111110001: M1r = 2'b01;
			14'b11010111110001: M1r = 2'b01;
			14'b00100111110001: M1r = 2'b00;
			14'b01100111110001: M1r = 2'b01;
			14'b10100111110001: M1r = 2'b01;
			14'b11100111110001: M1r = 2'b01;
			14'b00110111110001: M1r = 2'b00;
			14'b01110111110001: M1r = 2'b00;
			14'b10110111110001: M1r = 2'b00;
			14'b11110111110001: M1r = 2'b00;
			14'b00001011110001: M1r = 2'b10;
			14'b01001011110001: M1r = 2'b10;
			14'b10001011110001: M1r = 2'b10;
			14'b11001011110001: M1r = 2'b11;
			14'b00011011110001: M1r = 2'b10;
			14'b01011011110001: M1r = 2'b10;
			14'b10011011110001: M1r = 2'b10;
			14'b11011011110001: M1r = 2'b10;
			14'b00101011110001: M1r = 2'b01;
			14'b01101011110001: M1r = 2'b01;
			14'b10101011110001: M1r = 2'b01;
			14'b11101011110001: M1r = 2'b10;
			14'b00111011110001: M1r = 2'b01;
			14'b01111011110001: M1r = 2'b01;
			14'b10111011110001: M1r = 2'b01;
			14'b11111011110001: M1r = 2'b01;
			14'b00001111110001: M1r = 2'b11;
			14'b01001111110001: M1r = 2'b11;
			14'b10001111110001: M1r = 2'b11;
			14'b11001111110001: M1r = 2'b11;
			14'b00011111110001: M1r = 2'b10;
			14'b01011111110001: M1r = 2'b11;
			14'b10011111110001: M1r = 2'b11;
			14'b11011111110001: M1r = 2'b11;
			14'b00101111110001: M1r = 2'b10;
			14'b01101111110001: M1r = 2'b10;
			14'b10101111110001: M1r = 2'b10;
			14'b11101111110001: M1r = 2'b10;
			14'b00111111110001: M1r = 2'b01;
			14'b01111111110001: M1r = 2'b10;
			14'b10111111110001: M1r = 2'b10;
			14'b11111111110001: M1r = 2'b10;
			14'b00000000000101: M1r = 2'b00;
			14'b01000000000101: M1r = 2'b00;
			14'b10000000000101: M1r = 2'b00;
			14'b11000000000101: M1r = 2'b00;
			14'b00010000000101: M1r = 2'b00;
			14'b01010000000101: M1r = 2'b00;
			14'b10010000000101: M1r = 2'b00;
			14'b11010000000101: M1r = 2'b00;
			14'b00100000000101: M1r = 2'b00;
			14'b01100000000101: M1r = 2'b00;
			14'b10100000000101: M1r = 2'b00;
			14'b11100000000101: M1r = 2'b00;
			14'b00110000000101: M1r = 2'b00;
			14'b01110000000101: M1r = 2'b00;
			14'b10110000000101: M1r = 2'b00;
			14'b11110000000101: M1r = 2'b00;
			14'b00000100000101: M1r = 2'b00;
			14'b01000100000101: M1r = 2'b00;
			14'b10000100000101: M1r = 2'b00;
			14'b11000100000101: M1r = 2'b01;
			14'b00010100000101: M1r = 2'b00;
			14'b01010100000101: M1r = 2'b00;
			14'b10010100000101: M1r = 2'b00;
			14'b11010100000101: M1r = 2'b00;
			14'b00100100000101: M1r = 2'b00;
			14'b01100100000101: M1r = 2'b00;
			14'b10100100000101: M1r = 2'b00;
			14'b11100100000101: M1r = 2'b00;
			14'b00110100000101: M1r = 2'b00;
			14'b01110100000101: M1r = 2'b00;
			14'b10110100000101: M1r = 2'b00;
			14'b11110100000101: M1r = 2'b00;
			14'b00001000000101: M1r = 2'b01;
			14'b01001000000101: M1r = 2'b01;
			14'b10001000000101: M1r = 2'b01;
			14'b11001000000101: M1r = 2'b01;
			14'b00011000000101: M1r = 2'b00;
			14'b01011000000101: M1r = 2'b01;
			14'b10011000000101: M1r = 2'b01;
			14'b11011000000101: M1r = 2'b01;
			14'b00101000000101: M1r = 2'b00;
			14'b01101000000101: M1r = 2'b00;
			14'b10101000000101: M1r = 2'b00;
			14'b11101000000101: M1r = 2'b00;
			14'b00111000000101: M1r = 2'b00;
			14'b01111000000101: M1r = 2'b00;
			14'b10111000000101: M1r = 2'b00;
			14'b11111000000101: M1r = 2'b00;
			14'b00001100000101: M1r = 2'b10;
			14'b01001100000101: M1r = 2'b10;
			14'b10001100000101: M1r = 2'b10;
			14'b11001100000101: M1r = 2'b10;
			14'b00011100000101: M1r = 2'b01;
			14'b01011100000101: M1r = 2'b01;
			14'b10011100000101: M1r = 2'b01;
			14'b11011100000101: M1r = 2'b10;
			14'b00101100000101: M1r = 2'b01;
			14'b01101100000101: M1r = 2'b01;
			14'b10101100000101: M1r = 2'b01;
			14'b11101100000101: M1r = 2'b01;
			14'b00111100000101: M1r = 2'b00;
			14'b01111100000101: M1r = 2'b00;
			14'b10111100000101: M1r = 2'b00;
			14'b11111100000101: M1r = 2'b01;
			14'b00000001000101: M1r = 2'b00;
			14'b01000001000101: M1r = 2'b00;
			14'b10000001000101: M1r = 2'b00;
			14'b11000001000101: M1r = 2'b00;
			14'b00010001000101: M1r = 2'b00;
			14'b01010001000101: M1r = 2'b00;
			14'b10010001000101: M1r = 2'b00;
			14'b11010001000101: M1r = 2'b00;
			14'b00100001000101: M1r = 2'b00;
			14'b01100001000101: M1r = 2'b00;
			14'b10100001000101: M1r = 2'b00;
			14'b11100001000101: M1r = 2'b00;
			14'b00110001000101: M1r = 2'b00;
			14'b01110001000101: M1r = 2'b00;
			14'b10110001000101: M1r = 2'b00;
			14'b11110001000101: M1r = 2'b00;
			14'b00000101000101: M1r = 2'b00;
			14'b01000101000101: M1r = 2'b00;
			14'b10000101000101: M1r = 2'b00;
			14'b11000101000101: M1r = 2'b00;
			14'b00010101000101: M1r = 2'b00;
			14'b01010101000101: M1r = 2'b00;
			14'b10010101000101: M1r = 2'b00;
			14'b11010101000101: M1r = 2'b00;
			14'b00100101000101: M1r = 2'b00;
			14'b01100101000101: M1r = 2'b00;
			14'b10100101000101: M1r = 2'b00;
			14'b11100101000101: M1r = 2'b00;
			14'b00110101000101: M1r = 2'b00;
			14'b01110101000101: M1r = 2'b00;
			14'b10110101000101: M1r = 2'b00;
			14'b11110101000101: M1r = 2'b00;
			14'b00001001000101: M1r = 2'b01;
			14'b01001001000101: M1r = 2'b01;
			14'b10001001000101: M1r = 2'b01;
			14'b11001001000101: M1r = 2'b01;
			14'b00011001000101: M1r = 2'b00;
			14'b01011001000101: M1r = 2'b00;
			14'b10011001000101: M1r = 2'b00;
			14'b11011001000101: M1r = 2'b01;
			14'b00101001000101: M1r = 2'b00;
			14'b01101001000101: M1r = 2'b00;
			14'b10101001000101: M1r = 2'b00;
			14'b11101001000101: M1r = 2'b00;
			14'b00111001000101: M1r = 2'b00;
			14'b01111001000101: M1r = 2'b00;
			14'b10111001000101: M1r = 2'b00;
			14'b11111001000101: M1r = 2'b00;
			14'b00001101000101: M1r = 2'b01;
			14'b01001101000101: M1r = 2'b01;
			14'b10001101000101: M1r = 2'b10;
			14'b11001101000101: M1r = 2'b10;
			14'b00011101000101: M1r = 2'b01;
			14'b01011101000101: M1r = 2'b01;
			14'b10011101000101: M1r = 2'b01;
			14'b11011101000101: M1r = 2'b01;
			14'b00101101000101: M1r = 2'b00;
			14'b01101101000101: M1r = 2'b01;
			14'b10101101000101: M1r = 2'b01;
			14'b11101101000101: M1r = 2'b01;
			14'b00111101000101: M1r = 2'b00;
			14'b01111101000101: M1r = 2'b00;
			14'b10111101000101: M1r = 2'b00;
			14'b11111101000101: M1r = 2'b00;
			14'b00000010000101: M1r = 2'b00;
			14'b01000010000101: M1r = 2'b00;
			14'b10000010000101: M1r = 2'b00;
			14'b11000010000101: M1r = 2'b00;
			14'b00010010000101: M1r = 2'b00;
			14'b01010010000101: M1r = 2'b00;
			14'b10010010000101: M1r = 2'b00;
			14'b11010010000101: M1r = 2'b00;
			14'b00100010000101: M1r = 2'b00;
			14'b01100010000101: M1r = 2'b00;
			14'b10100010000101: M1r = 2'b00;
			14'b11100010000101: M1r = 2'b00;
			14'b00110010000101: M1r = 2'b00;
			14'b01110010000101: M1r = 2'b00;
			14'b10110010000101: M1r = 2'b00;
			14'b11110010000101: M1r = 2'b00;
			14'b00000110000101: M1r = 2'b00;
			14'b01000110000101: M1r = 2'b00;
			14'b10000110000101: M1r = 2'b00;
			14'b11000110000101: M1r = 2'b00;
			14'b00010110000101: M1r = 2'b00;
			14'b01010110000101: M1r = 2'b00;
			14'b10010110000101: M1r = 2'b00;
			14'b11010110000101: M1r = 2'b00;
			14'b00100110000101: M1r = 2'b00;
			14'b01100110000101: M1r = 2'b00;
			14'b10100110000101: M1r = 2'b00;
			14'b11100110000101: M1r = 2'b00;
			14'b00110110000101: M1r = 2'b00;
			14'b01110110000101: M1r = 2'b00;
			14'b10110110000101: M1r = 2'b00;
			14'b11110110000101: M1r = 2'b00;
			14'b00001010000101: M1r = 2'b00;
			14'b01001010000101: M1r = 2'b00;
			14'b10001010000101: M1r = 2'b01;
			14'b11001010000101: M1r = 2'b01;
			14'b00011010000101: M1r = 2'b00;
			14'b01011010000101: M1r = 2'b00;
			14'b10011010000101: M1r = 2'b00;
			14'b11011010000101: M1r = 2'b00;
			14'b00101010000101: M1r = 2'b00;
			14'b01101010000101: M1r = 2'b00;
			14'b10101010000101: M1r = 2'b00;
			14'b11101010000101: M1r = 2'b00;
			14'b00111010000101: M1r = 2'b00;
			14'b01111010000101: M1r = 2'b00;
			14'b10111010000101: M1r = 2'b00;
			14'b11111010000101: M1r = 2'b00;
			14'b00001110000101: M1r = 2'b01;
			14'b01001110000101: M1r = 2'b01;
			14'b10001110000101: M1r = 2'b01;
			14'b11001110000101: M1r = 2'b01;
			14'b00011110000101: M1r = 2'b01;
			14'b01011110000101: M1r = 2'b01;
			14'b10011110000101: M1r = 2'b01;
			14'b11011110000101: M1r = 2'b01;
			14'b00101110000101: M1r = 2'b00;
			14'b01101110000101: M1r = 2'b00;
			14'b10101110000101: M1r = 2'b00;
			14'b11101110000101: M1r = 2'b01;
			14'b00111110000101: M1r = 2'b00;
			14'b01111110000101: M1r = 2'b00;
			14'b10111110000101: M1r = 2'b00;
			14'b11111110000101: M1r = 2'b00;
			14'b00000011000101: M1r = 2'b00;
			14'b01000011000101: M1r = 2'b00;
			14'b10000011000101: M1r = 2'b00;
			14'b11000011000101: M1r = 2'b00;
			14'b00010011000101: M1r = 2'b00;
			14'b01010011000101: M1r = 2'b00;
			14'b10010011000101: M1r = 2'b00;
			14'b11010011000101: M1r = 2'b00;
			14'b00100011000101: M1r = 2'b00;
			14'b01100011000101: M1r = 2'b00;
			14'b10100011000101: M1r = 2'b00;
			14'b11100011000101: M1r = 2'b00;
			14'b00110011000101: M1r = 2'b00;
			14'b01110011000101: M1r = 2'b00;
			14'b10110011000101: M1r = 2'b00;
			14'b11110011000101: M1r = 2'b00;
			14'b00000111000101: M1r = 2'b00;
			14'b01000111000101: M1r = 2'b00;
			14'b10000111000101: M1r = 2'b00;
			14'b11000111000101: M1r = 2'b00;
			14'b00010111000101: M1r = 2'b00;
			14'b01010111000101: M1r = 2'b00;
			14'b10010111000101: M1r = 2'b00;
			14'b11010111000101: M1r = 2'b00;
			14'b00100111000101: M1r = 2'b00;
			14'b01100111000101: M1r = 2'b00;
			14'b10100111000101: M1r = 2'b00;
			14'b11100111000101: M1r = 2'b00;
			14'b00110111000101: M1r = 2'b00;
			14'b01110111000101: M1r = 2'b00;
			14'b10110111000101: M1r = 2'b00;
			14'b11110111000101: M1r = 2'b00;
			14'b00001011000101: M1r = 2'b00;
			14'b01001011000101: M1r = 2'b00;
			14'b10001011000101: M1r = 2'b00;
			14'b11001011000101: M1r = 2'b00;
			14'b00011011000101: M1r = 2'b00;
			14'b01011011000101: M1r = 2'b00;
			14'b10011011000101: M1r = 2'b00;
			14'b11011011000101: M1r = 2'b00;
			14'b00101011000101: M1r = 2'b00;
			14'b01101011000101: M1r = 2'b00;
			14'b10101011000101: M1r = 2'b00;
			14'b11101011000101: M1r = 2'b00;
			14'b00111011000101: M1r = 2'b00;
			14'b01111011000101: M1r = 2'b00;
			14'b10111011000101: M1r = 2'b00;
			14'b11111011000101: M1r = 2'b00;
			14'b00001111000101: M1r = 2'b01;
			14'b01001111000101: M1r = 2'b01;
			14'b10001111000101: M1r = 2'b01;
			14'b11001111000101: M1r = 2'b01;
			14'b00011111000101: M1r = 2'b00;
			14'b01011111000101: M1r = 2'b00;
			14'b10011111000101: M1r = 2'b01;
			14'b11011111000101: M1r = 2'b01;
			14'b00101111000101: M1r = 2'b00;
			14'b01101111000101: M1r = 2'b00;
			14'b10101111000101: M1r = 2'b00;
			14'b11101111000101: M1r = 2'b00;
			14'b00111111000101: M1r = 2'b00;
			14'b01111111000101: M1r = 2'b00;
			14'b10111111000101: M1r = 2'b00;
			14'b11111111000101: M1r = 2'b00;
			14'b00000000010101: M1r = 2'b00;
			14'b01000000010101: M1r = 2'b00;
			14'b10000000010101: M1r = 2'b00;
			14'b11000000010101: M1r = 2'b00;
			14'b00010000010101: M1r = 2'b00;
			14'b01010000010101: M1r = 2'b00;
			14'b10010000010101: M1r = 2'b00;
			14'b11010000010101: M1r = 2'b00;
			14'b00100000010101: M1r = 2'b00;
			14'b01100000010101: M1r = 2'b00;
			14'b10100000010101: M1r = 2'b00;
			14'b11100000010101: M1r = 2'b00;
			14'b00110000010101: M1r = 2'b00;
			14'b01110000010101: M1r = 2'b00;
			14'b10110000010101: M1r = 2'b00;
			14'b11110000010101: M1r = 2'b00;
			14'b00000100010101: M1r = 2'b01;
			14'b01000100010101: M1r = 2'b01;
			14'b10000100010101: M1r = 2'b01;
			14'b11000100010101: M1r = 2'b01;
			14'b00010100010101: M1r = 2'b00;
			14'b01010100010101: M1r = 2'b00;
			14'b10010100010101: M1r = 2'b00;
			14'b11010100010101: M1r = 2'b00;
			14'b00100100010101: M1r = 2'b00;
			14'b01100100010101: M1r = 2'b00;
			14'b10100100010101: M1r = 2'b00;
			14'b11100100010101: M1r = 2'b00;
			14'b00110100010101: M1r = 2'b00;
			14'b01110100010101: M1r = 2'b00;
			14'b10110100010101: M1r = 2'b00;
			14'b11110100010101: M1r = 2'b00;
			14'b00001000010101: M1r = 2'b01;
			14'b01001000010101: M1r = 2'b01;
			14'b10001000010101: M1r = 2'b10;
			14'b11001000010101: M1r = 2'b10;
			14'b00011000010101: M1r = 2'b01;
			14'b01011000010101: M1r = 2'b01;
			14'b10011000010101: M1r = 2'b01;
			14'b11011000010101: M1r = 2'b01;
			14'b00101000010101: M1r = 2'b00;
			14'b01101000010101: M1r = 2'b00;
			14'b10101000010101: M1r = 2'b01;
			14'b11101000010101: M1r = 2'b01;
			14'b00111000010101: M1r = 2'b00;
			14'b01111000010101: M1r = 2'b00;
			14'b10111000010101: M1r = 2'b00;
			14'b11111000010101: M1r = 2'b00;
			14'b00001100010101: M1r = 2'b10;
			14'b01001100010101: M1r = 2'b10;
			14'b10001100010101: M1r = 2'b10;
			14'b11001100010101: M1r = 2'b10;
			14'b00011100010101: M1r = 2'b10;
			14'b01011100010101: M1r = 2'b10;
			14'b10011100010101: M1r = 2'b10;
			14'b11011100010101: M1r = 2'b10;
			14'b00101100010101: M1r = 2'b01;
			14'b01101100010101: M1r = 2'b01;
			14'b10101100010101: M1r = 2'b01;
			14'b11101100010101: M1r = 2'b10;
			14'b00111100010101: M1r = 2'b01;
			14'b01111100010101: M1r = 2'b01;
			14'b10111100010101: M1r = 2'b01;
			14'b11111100010101: M1r = 2'b01;
			14'b00000001010101: M1r = 2'b00;
			14'b01000001010101: M1r = 2'b00;
			14'b10000001010101: M1r = 2'b00;
			14'b11000001010101: M1r = 2'b00;
			14'b00010001010101: M1r = 2'b00;
			14'b01010001010101: M1r = 2'b00;
			14'b10010001010101: M1r = 2'b00;
			14'b11010001010101: M1r = 2'b00;
			14'b00100001010101: M1r = 2'b00;
			14'b01100001010101: M1r = 2'b00;
			14'b10100001010101: M1r = 2'b00;
			14'b11100001010101: M1r = 2'b00;
			14'b00110001010101: M1r = 2'b00;
			14'b01110001010101: M1r = 2'b00;
			14'b10110001010101: M1r = 2'b00;
			14'b11110001010101: M1r = 2'b00;
			14'b00000101010101: M1r = 2'b00;
			14'b01000101010101: M1r = 2'b00;
			14'b10000101010101: M1r = 2'b01;
			14'b11000101010101: M1r = 2'b01;
			14'b00010101010101: M1r = 2'b00;
			14'b01010101010101: M1r = 2'b00;
			14'b10010101010101: M1r = 2'b00;
			14'b11010101010101: M1r = 2'b00;
			14'b00100101010101: M1r = 2'b00;
			14'b01100101010101: M1r = 2'b00;
			14'b10100101010101: M1r = 2'b00;
			14'b11100101010101: M1r = 2'b00;
			14'b00110101010101: M1r = 2'b00;
			14'b01110101010101: M1r = 2'b00;
			14'b10110101010101: M1r = 2'b00;
			14'b11110101010101: M1r = 2'b00;
			14'b00001001010101: M1r = 2'b01;
			14'b01001001010101: M1r = 2'b01;
			14'b10001001010101: M1r = 2'b01;
			14'b11001001010101: M1r = 2'b01;
			14'b00011001010101: M1r = 2'b01;
			14'b01011001010101: M1r = 2'b01;
			14'b10011001010101: M1r = 2'b01;
			14'b11011001010101: M1r = 2'b01;
			14'b00101001010101: M1r = 2'b00;
			14'b01101001010101: M1r = 2'b00;
			14'b10101001010101: M1r = 2'b00;
			14'b11101001010101: M1r = 2'b00;
			14'b00111001010101: M1r = 2'b00;
			14'b01111001010101: M1r = 2'b00;
			14'b10111001010101: M1r = 2'b00;
			14'b11111001010101: M1r = 2'b00;
			14'b00001101010101: M1r = 2'b10;
			14'b01001101010101: M1r = 2'b10;
			14'b10001101010101: M1r = 2'b10;
			14'b11001101010101: M1r = 2'b10;
			14'b00011101010101: M1r = 2'b01;
			14'b01011101010101: M1r = 2'b01;
			14'b10011101010101: M1r = 2'b10;
			14'b11011101010101: M1r = 2'b10;
			14'b00101101010101: M1r = 2'b01;
			14'b01101101010101: M1r = 2'b01;
			14'b10101101010101: M1r = 2'b01;
			14'b11101101010101: M1r = 2'b01;
			14'b00111101010101: M1r = 2'b00;
			14'b01111101010101: M1r = 2'b00;
			14'b10111101010101: M1r = 2'b01;
			14'b11111101010101: M1r = 2'b01;
			14'b00000010010101: M1r = 2'b00;
			14'b01000010010101: M1r = 2'b00;
			14'b10000010010101: M1r = 2'b00;
			14'b11000010010101: M1r = 2'b00;
			14'b00010010010101: M1r = 2'b00;
			14'b01010010010101: M1r = 2'b00;
			14'b10010010010101: M1r = 2'b00;
			14'b11010010010101: M1r = 2'b00;
			14'b00100010010101: M1r = 2'b00;
			14'b01100010010101: M1r = 2'b00;
			14'b10100010010101: M1r = 2'b00;
			14'b11100010010101: M1r = 2'b00;
			14'b00110010010101: M1r = 2'b00;
			14'b01110010010101: M1r = 2'b00;
			14'b10110010010101: M1r = 2'b00;
			14'b11110010010101: M1r = 2'b00;
			14'b00000110010101: M1r = 2'b00;
			14'b01000110010101: M1r = 2'b00;
			14'b10000110010101: M1r = 2'b00;
			14'b11000110010101: M1r = 2'b00;
			14'b00010110010101: M1r = 2'b00;
			14'b01010110010101: M1r = 2'b00;
			14'b10010110010101: M1r = 2'b00;
			14'b11010110010101: M1r = 2'b00;
			14'b00100110010101: M1r = 2'b00;
			14'b01100110010101: M1r = 2'b00;
			14'b10100110010101: M1r = 2'b00;
			14'b11100110010101: M1r = 2'b00;
			14'b00110110010101: M1r = 2'b00;
			14'b01110110010101: M1r = 2'b00;
			14'b10110110010101: M1r = 2'b00;
			14'b11110110010101: M1r = 2'b00;
			14'b00001010010101: M1r = 2'b01;
			14'b01001010010101: M1r = 2'b01;
			14'b10001010010101: M1r = 2'b01;
			14'b11001010010101: M1r = 2'b01;
			14'b00011010010101: M1r = 2'b00;
			14'b01011010010101: M1r = 2'b00;
			14'b10011010010101: M1r = 2'b01;
			14'b11011010010101: M1r = 2'b01;
			14'b00101010010101: M1r = 2'b00;
			14'b01101010010101: M1r = 2'b00;
			14'b10101010010101: M1r = 2'b00;
			14'b11101010010101: M1r = 2'b00;
			14'b00111010010101: M1r = 2'b00;
			14'b01111010010101: M1r = 2'b00;
			14'b10111010010101: M1r = 2'b00;
			14'b11111010010101: M1r = 2'b00;
			14'b00001110010101: M1r = 2'b01;
			14'b01001110010101: M1r = 2'b10;
			14'b10001110010101: M1r = 2'b10;
			14'b11001110010101: M1r = 2'b10;
			14'b00011110010101: M1r = 2'b01;
			14'b01011110010101: M1r = 2'b01;
			14'b10011110010101: M1r = 2'b01;
			14'b11011110010101: M1r = 2'b01;
			14'b00101110010101: M1r = 2'b01;
			14'b01101110010101: M1r = 2'b01;
			14'b10101110010101: M1r = 2'b01;
			14'b11101110010101: M1r = 2'b01;
			14'b00111110010101: M1r = 2'b00;
			14'b01111110010101: M1r = 2'b00;
			14'b10111110010101: M1r = 2'b00;
			14'b11111110010101: M1r = 2'b00;
			14'b00000011010101: M1r = 2'b00;
			14'b01000011010101: M1r = 2'b00;
			14'b10000011010101: M1r = 2'b00;
			14'b11000011010101: M1r = 2'b00;
			14'b00010011010101: M1r = 2'b00;
			14'b01010011010101: M1r = 2'b00;
			14'b10010011010101: M1r = 2'b00;
			14'b11010011010101: M1r = 2'b00;
			14'b00100011010101: M1r = 2'b00;
			14'b01100011010101: M1r = 2'b00;
			14'b10100011010101: M1r = 2'b00;
			14'b11100011010101: M1r = 2'b00;
			14'b00110011010101: M1r = 2'b00;
			14'b01110011010101: M1r = 2'b00;
			14'b10110011010101: M1r = 2'b00;
			14'b11110011010101: M1r = 2'b00;
			14'b00000111010101: M1r = 2'b00;
			14'b01000111010101: M1r = 2'b00;
			14'b10000111010101: M1r = 2'b00;
			14'b11000111010101: M1r = 2'b00;
			14'b00010111010101: M1r = 2'b00;
			14'b01010111010101: M1r = 2'b00;
			14'b10010111010101: M1r = 2'b00;
			14'b11010111010101: M1r = 2'b00;
			14'b00100111010101: M1r = 2'b00;
			14'b01100111010101: M1r = 2'b00;
			14'b10100111010101: M1r = 2'b00;
			14'b11100111010101: M1r = 2'b00;
			14'b00110111010101: M1r = 2'b00;
			14'b01110111010101: M1r = 2'b00;
			14'b10110111010101: M1r = 2'b00;
			14'b11110111010101: M1r = 2'b00;
			14'b00001011010101: M1r = 2'b00;
			14'b01001011010101: M1r = 2'b01;
			14'b10001011010101: M1r = 2'b01;
			14'b11001011010101: M1r = 2'b01;
			14'b00011011010101: M1r = 2'b00;
			14'b01011011010101: M1r = 2'b00;
			14'b10011011010101: M1r = 2'b00;
			14'b11011011010101: M1r = 2'b00;
			14'b00101011010101: M1r = 2'b00;
			14'b01101011010101: M1r = 2'b00;
			14'b10101011010101: M1r = 2'b00;
			14'b11101011010101: M1r = 2'b00;
			14'b00111011010101: M1r = 2'b00;
			14'b01111011010101: M1r = 2'b00;
			14'b10111011010101: M1r = 2'b00;
			14'b11111011010101: M1r = 2'b00;
			14'b00001111010101: M1r = 2'b01;
			14'b01001111010101: M1r = 2'b01;
			14'b10001111010101: M1r = 2'b01;
			14'b11001111010101: M1r = 2'b10;
			14'b00011111010101: M1r = 2'b01;
			14'b01011111010101: M1r = 2'b01;
			14'b10011111010101: M1r = 2'b01;
			14'b11011111010101: M1r = 2'b01;
			14'b00101111010101: M1r = 2'b00;
			14'b01101111010101: M1r = 2'b00;
			14'b10101111010101: M1r = 2'b01;
			14'b11101111010101: M1r = 2'b01;
			14'b00111111010101: M1r = 2'b00;
			14'b01111111010101: M1r = 2'b00;
			14'b10111111010101: M1r = 2'b00;
			14'b11111111010101: M1r = 2'b00;
			14'b00000000100101: M1r = 2'b00;
			14'b01000000100101: M1r = 2'b00;
			14'b10000000100101: M1r = 2'b00;
			14'b11000000100101: M1r = 2'b01;
			14'b00010000100101: M1r = 2'b00;
			14'b01010000100101: M1r = 2'b00;
			14'b10010000100101: M1r = 2'b00;
			14'b11010000100101: M1r = 2'b00;
			14'b00100000100101: M1r = 2'b00;
			14'b01100000100101: M1r = 2'b00;
			14'b10100000100101: M1r = 2'b00;
			14'b11100000100101: M1r = 2'b00;
			14'b00110000100101: M1r = 2'b00;
			14'b01110000100101: M1r = 2'b00;
			14'b10110000100101: M1r = 2'b00;
			14'b11110000100101: M1r = 2'b00;
			14'b00000100100101: M1r = 2'b01;
			14'b01000100100101: M1r = 2'b01;
			14'b10000100100101: M1r = 2'b01;
			14'b11000100100101: M1r = 2'b01;
			14'b00010100100101: M1r = 2'b00;
			14'b01010100100101: M1r = 2'b01;
			14'b10010100100101: M1r = 2'b01;
			14'b11010100100101: M1r = 2'b01;
			14'b00100100100101: M1r = 2'b00;
			14'b01100100100101: M1r = 2'b00;
			14'b10100100100101: M1r = 2'b00;
			14'b11100100100101: M1r = 2'b00;
			14'b00110100100101: M1r = 2'b00;
			14'b01110100100101: M1r = 2'b00;
			14'b10110100100101: M1r = 2'b00;
			14'b11110100100101: M1r = 2'b00;
			14'b00001000100101: M1r = 2'b10;
			14'b01001000100101: M1r = 2'b10;
			14'b10001000100101: M1r = 2'b10;
			14'b11001000100101: M1r = 2'b10;
			14'b00011000100101: M1r = 2'b01;
			14'b01011000100101: M1r = 2'b01;
			14'b10011000100101: M1r = 2'b10;
			14'b11011000100101: M1r = 2'b10;
			14'b00101000100101: M1r = 2'b01;
			14'b01101000100101: M1r = 2'b01;
			14'b10101000100101: M1r = 2'b01;
			14'b11101000100101: M1r = 2'b01;
			14'b00111000100101: M1r = 2'b00;
			14'b01111000100101: M1r = 2'b00;
			14'b10111000100101: M1r = 2'b01;
			14'b11111000100101: M1r = 2'b01;
			14'b00001100100101: M1r = 2'b10;
			14'b01001100100101: M1r = 2'b11;
			14'b10001100100101: M1r = 2'b11;
			14'b11001100100101: M1r = 2'b11;
			14'b00011100100101: M1r = 2'b10;
			14'b01011100100101: M1r = 2'b10;
			14'b10011100100101: M1r = 2'b10;
			14'b11011100100101: M1r = 2'b10;
			14'b00101100100101: M1r = 2'b01;
			14'b01101100100101: M1r = 2'b10;
			14'b10101100100101: M1r = 2'b10;
			14'b11101100100101: M1r = 2'b10;
			14'b00111100100101: M1r = 2'b01;
			14'b01111100100101: M1r = 2'b01;
			14'b10111100100101: M1r = 2'b01;
			14'b11111100100101: M1r = 2'b01;
			14'b00000001100101: M1r = 2'b00;
			14'b01000001100101: M1r = 2'b00;
			14'b10000001100101: M1r = 2'b00;
			14'b11000001100101: M1r = 2'b00;
			14'b00010001100101: M1r = 2'b00;
			14'b01010001100101: M1r = 2'b00;
			14'b10010001100101: M1r = 2'b00;
			14'b11010001100101: M1r = 2'b00;
			14'b00100001100101: M1r = 2'b00;
			14'b01100001100101: M1r = 2'b00;
			14'b10100001100101: M1r = 2'b00;
			14'b11100001100101: M1r = 2'b00;
			14'b00110001100101: M1r = 2'b00;
			14'b01110001100101: M1r = 2'b00;
			14'b10110001100101: M1r = 2'b00;
			14'b11110001100101: M1r = 2'b00;
			14'b00000101100101: M1r = 2'b01;
			14'b01000101100101: M1r = 2'b01;
			14'b10000101100101: M1r = 2'b01;
			14'b11000101100101: M1r = 2'b01;
			14'b00010101100101: M1r = 2'b00;
			14'b01010101100101: M1r = 2'b00;
			14'b10010101100101: M1r = 2'b00;
			14'b11010101100101: M1r = 2'b01;
			14'b00100101100101: M1r = 2'b00;
			14'b01100101100101: M1r = 2'b00;
			14'b10100101100101: M1r = 2'b00;
			14'b11100101100101: M1r = 2'b00;
			14'b00110101100101: M1r = 2'b00;
			14'b01110101100101: M1r = 2'b00;
			14'b10110101100101: M1r = 2'b00;
			14'b11110101100101: M1r = 2'b00;
			14'b00001001100101: M1r = 2'b01;
			14'b01001001100101: M1r = 2'b10;
			14'b10001001100101: M1r = 2'b10;
			14'b11001001100101: M1r = 2'b10;
			14'b00011001100101: M1r = 2'b01;
			14'b01011001100101: M1r = 2'b01;
			14'b10011001100101: M1r = 2'b01;
			14'b11011001100101: M1r = 2'b01;
			14'b00101001100101: M1r = 2'b00;
			14'b01101001100101: M1r = 2'b01;
			14'b10101001100101: M1r = 2'b01;
			14'b11101001100101: M1r = 2'b01;
			14'b00111001100101: M1r = 2'b00;
			14'b01111001100101: M1r = 2'b00;
			14'b10111001100101: M1r = 2'b00;
			14'b11111001100101: M1r = 2'b00;
			14'b00001101100101: M1r = 2'b10;
			14'b01001101100101: M1r = 2'b10;
			14'b10001101100101: M1r = 2'b10;
			14'b11001101100101: M1r = 2'b11;
			14'b00011101100101: M1r = 2'b10;
			14'b01011101100101: M1r = 2'b10;
			14'b10011101100101: M1r = 2'b10;
			14'b11011101100101: M1r = 2'b10;
			14'b00101101100101: M1r = 2'b01;
			14'b01101101100101: M1r = 2'b01;
			14'b10101101100101: M1r = 2'b10;
			14'b11101101100101: M1r = 2'b10;
			14'b00111101100101: M1r = 2'b01;
			14'b01111101100101: M1r = 2'b01;
			14'b10111101100101: M1r = 2'b01;
			14'b11111101100101: M1r = 2'b01;
			14'b00000010100101: M1r = 2'b00;
			14'b01000010100101: M1r = 2'b00;
			14'b10000010100101: M1r = 2'b00;
			14'b11000010100101: M1r = 2'b00;
			14'b00010010100101: M1r = 2'b00;
			14'b01010010100101: M1r = 2'b00;
			14'b10010010100101: M1r = 2'b00;
			14'b11010010100101: M1r = 2'b00;
			14'b00100010100101: M1r = 2'b00;
			14'b01100010100101: M1r = 2'b00;
			14'b10100010100101: M1r = 2'b00;
			14'b11100010100101: M1r = 2'b00;
			14'b00110010100101: M1r = 2'b00;
			14'b01110010100101: M1r = 2'b00;
			14'b10110010100101: M1r = 2'b00;
			14'b11110010100101: M1r = 2'b00;
			14'b00000110100101: M1r = 2'b00;
			14'b01000110100101: M1r = 2'b01;
			14'b10000110100101: M1r = 2'b01;
			14'b11000110100101: M1r = 2'b01;
			14'b00010110100101: M1r = 2'b00;
			14'b01010110100101: M1r = 2'b00;
			14'b10010110100101: M1r = 2'b00;
			14'b11010110100101: M1r = 2'b00;
			14'b00100110100101: M1r = 2'b00;
			14'b01100110100101: M1r = 2'b00;
			14'b10100110100101: M1r = 2'b00;
			14'b11100110100101: M1r = 2'b00;
			14'b00110110100101: M1r = 2'b00;
			14'b01110110100101: M1r = 2'b00;
			14'b10110110100101: M1r = 2'b00;
			14'b11110110100101: M1r = 2'b00;
			14'b00001010100101: M1r = 2'b01;
			14'b01001010100101: M1r = 2'b01;
			14'b10001010100101: M1r = 2'b01;
			14'b11001010100101: M1r = 2'b10;
			14'b00011010100101: M1r = 2'b01;
			14'b01011010100101: M1r = 2'b01;
			14'b10011010100101: M1r = 2'b01;
			14'b11011010100101: M1r = 2'b01;
			14'b00101010100101: M1r = 2'b00;
			14'b01101010100101: M1r = 2'b00;
			14'b10101010100101: M1r = 2'b01;
			14'b11101010100101: M1r = 2'b01;
			14'b00111010100101: M1r = 2'b00;
			14'b01111010100101: M1r = 2'b00;
			14'b10111010100101: M1r = 2'b00;
			14'b11111010100101: M1r = 2'b00;
			14'b00001110100101: M1r = 2'b10;
			14'b01001110100101: M1r = 2'b10;
			14'b10001110100101: M1r = 2'b10;
			14'b11001110100101: M1r = 2'b10;
			14'b00011110100101: M1r = 2'b01;
			14'b01011110100101: M1r = 2'b10;
			14'b10011110100101: M1r = 2'b10;
			14'b11011110100101: M1r = 2'b10;
			14'b00101110100101: M1r = 2'b01;
			14'b01101110100101: M1r = 2'b01;
			14'b10101110100101: M1r = 2'b01;
			14'b11101110100101: M1r = 2'b01;
			14'b00111110100101: M1r = 2'b00;
			14'b01111110100101: M1r = 2'b01;
			14'b10111110100101: M1r = 2'b01;
			14'b11111110100101: M1r = 2'b01;
			14'b00000011100101: M1r = 2'b00;
			14'b01000011100101: M1r = 2'b00;
			14'b10000011100101: M1r = 2'b00;
			14'b11000011100101: M1r = 2'b00;
			14'b00010011100101: M1r = 2'b00;
			14'b01010011100101: M1r = 2'b00;
			14'b10010011100101: M1r = 2'b00;
			14'b11010011100101: M1r = 2'b00;
			14'b00100011100101: M1r = 2'b00;
			14'b01100011100101: M1r = 2'b00;
			14'b10100011100101: M1r = 2'b00;
			14'b11100011100101: M1r = 2'b00;
			14'b00110011100101: M1r = 2'b00;
			14'b01110011100101: M1r = 2'b00;
			14'b10110011100101: M1r = 2'b00;
			14'b11110011100101: M1r = 2'b00;
			14'b00000111100101: M1r = 2'b00;
			14'b01000111100101: M1r = 2'b00;
			14'b10000111100101: M1r = 2'b00;
			14'b11000111100101: M1r = 2'b01;
			14'b00010111100101: M1r = 2'b00;
			14'b01010111100101: M1r = 2'b00;
			14'b10010111100101: M1r = 2'b00;
			14'b11010111100101: M1r = 2'b00;
			14'b00100111100101: M1r = 2'b00;
			14'b01100111100101: M1r = 2'b00;
			14'b10100111100101: M1r = 2'b00;
			14'b11100111100101: M1r = 2'b00;
			14'b00110111100101: M1r = 2'b00;
			14'b01110111100101: M1r = 2'b00;
			14'b10110111100101: M1r = 2'b00;
			14'b11110111100101: M1r = 2'b00;
			14'b00001011100101: M1r = 2'b01;
			14'b01001011100101: M1r = 2'b01;
			14'b10001011100101: M1r = 2'b01;
			14'b11001011100101: M1r = 2'b01;
			14'b00011011100101: M1r = 2'b00;
			14'b01011011100101: M1r = 2'b01;
			14'b10011011100101: M1r = 2'b01;
			14'b11011011100101: M1r = 2'b01;
			14'b00101011100101: M1r = 2'b00;
			14'b01101011100101: M1r = 2'b00;
			14'b10101011100101: M1r = 2'b00;
			14'b11101011100101: M1r = 2'b00;
			14'b00111011100101: M1r = 2'b00;
			14'b01111011100101: M1r = 2'b00;
			14'b10111011100101: M1r = 2'b00;
			14'b11111011100101: M1r = 2'b00;
			14'b00001111100101: M1r = 2'b10;
			14'b01001111100101: M1r = 2'b10;
			14'b10001111100101: M1r = 2'b10;
			14'b11001111100101: M1r = 2'b10;
			14'b00011111100101: M1r = 2'b01;
			14'b01011111100101: M1r = 2'b01;
			14'b10011111100101: M1r = 2'b01;
			14'b11011111100101: M1r = 2'b10;
			14'b00101111100101: M1r = 2'b01;
			14'b01101111100101: M1r = 2'b01;
			14'b10101111100101: M1r = 2'b01;
			14'b11101111100101: M1r = 2'b01;
			14'b00111111100101: M1r = 2'b00;
			14'b01111111100101: M1r = 2'b00;
			14'b10111111100101: M1r = 2'b01;
			14'b11111111100101: M1r = 2'b01;
			14'b00000000110101: M1r = 2'b01;
			14'b01000000110101: M1r = 2'b01;
			14'b10000000110101: M1r = 2'b01;
			14'b11000000110101: M1r = 2'b01;
			14'b00010000110101: M1r = 2'b00;
			14'b01010000110101: M1r = 2'b00;
			14'b10010000110101: M1r = 2'b00;
			14'b11010000110101: M1r = 2'b01;
			14'b00100000110101: M1r = 2'b00;
			14'b01100000110101: M1r = 2'b00;
			14'b10100000110101: M1r = 2'b00;
			14'b11100000110101: M1r = 2'b00;
			14'b00110000110101: M1r = 2'b00;
			14'b01110000110101: M1r = 2'b00;
			14'b10110000110101: M1r = 2'b00;
			14'b11110000110101: M1r = 2'b00;
			14'b00000100110101: M1r = 2'b01;
			14'b01000100110101: M1r = 2'b10;
			14'b10000100110101: M1r = 2'b10;
			14'b11000100110101: M1r = 2'b10;
			14'b00010100110101: M1r = 2'b01;
			14'b01010100110101: M1r = 2'b01;
			14'b10010100110101: M1r = 2'b01;
			14'b11010100110101: M1r = 2'b01;
			14'b00100100110101: M1r = 2'b00;
			14'b01100100110101: M1r = 2'b01;
			14'b10100100110101: M1r = 2'b01;
			14'b11100100110101: M1r = 2'b01;
			14'b00110100110101: M1r = 2'b00;
			14'b01110100110101: M1r = 2'b00;
			14'b10110100110101: M1r = 2'b00;
			14'b11110100110101: M1r = 2'b00;
			14'b00001000110101: M1r = 2'b10;
			14'b01001000110101: M1r = 2'b10;
			14'b10001000110101: M1r = 2'b10;
			14'b11001000110101: M1r = 2'b11;
			14'b00011000110101: M1r = 2'b10;
			14'b01011000110101: M1r = 2'b10;
			14'b10011000110101: M1r = 2'b10;
			14'b11011000110101: M1r = 2'b10;
			14'b00101000110101: M1r = 2'b01;
			14'b01101000110101: M1r = 2'b01;
			14'b10101000110101: M1r = 2'b01;
			14'b11101000110101: M1r = 2'b10;
			14'b00111000110101: M1r = 2'b01;
			14'b01111000110101: M1r = 2'b01;
			14'b10111000110101: M1r = 2'b01;
			14'b11111000110101: M1r = 2'b01;
			14'b00001100110101: M1r = 2'b11;
			14'b01001100110101: M1r = 2'b11;
			14'b10001100110101: M1r = 2'b11;
			14'b11001100110101: M1r = 2'b11;
			14'b00011100110101: M1r = 2'b10;
			14'b01011100110101: M1r = 2'b11;
			14'b10011100110101: M1r = 2'b11;
			14'b11011100110101: M1r = 2'b11;
			14'b00101100110101: M1r = 2'b10;
			14'b01101100110101: M1r = 2'b10;
			14'b10101100110101: M1r = 2'b10;
			14'b11101100110101: M1r = 2'b10;
			14'b00111100110101: M1r = 2'b01;
			14'b01111100110101: M1r = 2'b10;
			14'b10111100110101: M1r = 2'b10;
			14'b11111100110101: M1r = 2'b10;
			14'b00000001110101: M1r = 2'b00;
			14'b01000001110101: M1r = 2'b01;
			14'b10000001110101: M1r = 2'b01;
			14'b11000001110101: M1r = 2'b01;
			14'b00010001110101: M1r = 2'b00;
			14'b01010001110101: M1r = 2'b00;
			14'b10010001110101: M1r = 2'b00;
			14'b11010001110101: M1r = 2'b00;
			14'b00100001110101: M1r = 2'b00;
			14'b01100001110101: M1r = 2'b00;
			14'b10100001110101: M1r = 2'b00;
			14'b11100001110101: M1r = 2'b00;
			14'b00110001110101: M1r = 2'b00;
			14'b01110001110101: M1r = 2'b00;
			14'b10110001110101: M1r = 2'b00;
			14'b11110001110101: M1r = 2'b00;
			14'b00000101110101: M1r = 2'b01;
			14'b01000101110101: M1r = 2'b01;
			14'b10000101110101: M1r = 2'b01;
			14'b11000101110101: M1r = 2'b10;
			14'b00010101110101: M1r = 2'b01;
			14'b01010101110101: M1r = 2'b01;
			14'b10010101110101: M1r = 2'b01;
			14'b11010101110101: M1r = 2'b01;
			14'b00100101110101: M1r = 2'b00;
			14'b01100101110101: M1r = 2'b00;
			14'b10100101110101: M1r = 2'b00;
			14'b11100101110101: M1r = 2'b01;
			14'b00110101110101: M1r = 2'b00;
			14'b01110101110101: M1r = 2'b00;
			14'b10110101110101: M1r = 2'b00;
			14'b11110101110101: M1r = 2'b00;
			14'b00001001110101: M1r = 2'b10;
			14'b01001001110101: M1r = 2'b10;
			14'b10001001110101: M1r = 2'b10;
			14'b11001001110101: M1r = 2'b10;
			14'b00011001110101: M1r = 2'b01;
			14'b01011001110101: M1r = 2'b10;
			14'b10011001110101: M1r = 2'b10;
			14'b11011001110101: M1r = 2'b10;
			14'b00101001110101: M1r = 2'b01;
			14'b01101001110101: M1r = 2'b01;
			14'b10101001110101: M1r = 2'b01;
			14'b11101001110101: M1r = 2'b01;
			14'b00111001110101: M1r = 2'b00;
			14'b01111001110101: M1r = 2'b01;
			14'b10111001110101: M1r = 2'b01;
			14'b11111001110101: M1r = 2'b01;
			14'b00001101110101: M1r = 2'b11;
			14'b01001101110101: M1r = 2'b11;
			14'b10001101110101: M1r = 2'b11;
			14'b11001101110101: M1r = 2'b11;
			14'b00011101110101: M1r = 2'b10;
			14'b01011101110101: M1r = 2'b10;
			14'b10011101110101: M1r = 2'b10;
			14'b11011101110101: M1r = 2'b11;
			14'b00101101110101: M1r = 2'b10;
			14'b01101101110101: M1r = 2'b10;
			14'b10101101110101: M1r = 2'b10;
			14'b11101101110101: M1r = 2'b10;
			14'b00111101110101: M1r = 2'b01;
			14'b01111101110101: M1r = 2'b01;
			14'b10111101110101: M1r = 2'b01;
			14'b11111101110101: M1r = 2'b10;
			14'b00000010110101: M1r = 2'b00;
			14'b01000010110101: M1r = 2'b00;
			14'b10000010110101: M1r = 2'b00;
			14'b11000010110101: M1r = 2'b01;
			14'b00010010110101: M1r = 2'b00;
			14'b01010010110101: M1r = 2'b00;
			14'b10010010110101: M1r = 2'b00;
			14'b11010010110101: M1r = 2'b00;
			14'b00100010110101: M1r = 2'b00;
			14'b01100010110101: M1r = 2'b00;
			14'b10100010110101: M1r = 2'b00;
			14'b11100010110101: M1r = 2'b00;
			14'b00110010110101: M1r = 2'b00;
			14'b01110010110101: M1r = 2'b00;
			14'b10110010110101: M1r = 2'b00;
			14'b11110010110101: M1r = 2'b00;
			14'b00000110110101: M1r = 2'b01;
			14'b01000110110101: M1r = 2'b01;
			14'b10000110110101: M1r = 2'b01;
			14'b11000110110101: M1r = 2'b01;
			14'b00010110110101: M1r = 2'b00;
			14'b01010110110101: M1r = 2'b01;
			14'b10010110110101: M1r = 2'b01;
			14'b11010110110101: M1r = 2'b01;
			14'b00100110110101: M1r = 2'b00;
			14'b01100110110101: M1r = 2'b00;
			14'b10100110110101: M1r = 2'b00;
			14'b11100110110101: M1r = 2'b00;
			14'b00110110110101: M1r = 2'b00;
			14'b01110110110101: M1r = 2'b00;
			14'b10110110110101: M1r = 2'b00;
			14'b11110110110101: M1r = 2'b00;
			14'b00001010110101: M1r = 2'b10;
			14'b01001010110101: M1r = 2'b10;
			14'b10001010110101: M1r = 2'b10;
			14'b11001010110101: M1r = 2'b10;
			14'b00011010110101: M1r = 2'b01;
			14'b01011010110101: M1r = 2'b01;
			14'b10011010110101: M1r = 2'b01;
			14'b11011010110101: M1r = 2'b10;
			14'b00101010110101: M1r = 2'b01;
			14'b01101010110101: M1r = 2'b01;
			14'b10101010110101: M1r = 2'b01;
			14'b11101010110101: M1r = 2'b01;
			14'b00111010110101: M1r = 2'b00;
			14'b01111010110101: M1r = 2'b00;
			14'b10111010110101: M1r = 2'b00;
			14'b11111010110101: M1r = 2'b01;
			14'b00001110110101: M1r = 2'b10;
			14'b01001110110101: M1r = 2'b10;
			14'b10001110110101: M1r = 2'b11;
			14'b11001110110101: M1r = 2'b11;
			14'b00011110110101: M1r = 2'b10;
			14'b01011110110101: M1r = 2'b10;
			14'b10011110110101: M1r = 2'b10;
			14'b11011110110101: M1r = 2'b10;
			14'b00101110110101: M1r = 2'b01;
			14'b01101110110101: M1r = 2'b10;
			14'b10101110110101: M1r = 2'b10;
			14'b11101110110101: M1r = 2'b10;
			14'b00111110110101: M1r = 2'b01;
			14'b01111110110101: M1r = 2'b01;
			14'b10111110110101: M1r = 2'b01;
			14'b11111110110101: M1r = 2'b01;
			14'b00000011110101: M1r = 2'b00;
			14'b01000011110101: M1r = 2'b00;
			14'b10000011110101: M1r = 2'b00;
			14'b11000011110101: M1r = 2'b00;
			14'b00010011110101: M1r = 2'b00;
			14'b01010011110101: M1r = 2'b00;
			14'b10010011110101: M1r = 2'b00;
			14'b11010011110101: M1r = 2'b00;
			14'b00100011110101: M1r = 2'b00;
			14'b01100011110101: M1r = 2'b00;
			14'b10100011110101: M1r = 2'b00;
			14'b11100011110101: M1r = 2'b00;
			14'b00110011110101: M1r = 2'b00;
			14'b01110011110101: M1r = 2'b00;
			14'b10110011110101: M1r = 2'b00;
			14'b11110011110101: M1r = 2'b00;
			14'b00000111110101: M1r = 2'b01;
			14'b01000111110101: M1r = 2'b01;
			14'b10000111110101: M1r = 2'b01;
			14'b11000111110101: M1r = 2'b01;
			14'b00010111110101: M1r = 2'b00;
			14'b01010111110101: M1r = 2'b00;
			14'b10010111110101: M1r = 2'b00;
			14'b11010111110101: M1r = 2'b01;
			14'b00100111110101: M1r = 2'b00;
			14'b01100111110101: M1r = 2'b00;
			14'b10100111110101: M1r = 2'b00;
			14'b11100111110101: M1r = 2'b00;
			14'b00110111110101: M1r = 2'b00;
			14'b01110111110101: M1r = 2'b00;
			14'b10110111110101: M1r = 2'b00;
			14'b11110111110101: M1r = 2'b00;
			14'b00001011110101: M1r = 2'b01;
			14'b01001011110101: M1r = 2'b01;
			14'b10001011110101: M1r = 2'b10;
			14'b11001011110101: M1r = 2'b10;
			14'b00011011110101: M1r = 2'b01;
			14'b01011011110101: M1r = 2'b01;
			14'b10011011110101: M1r = 2'b01;
			14'b11011011110101: M1r = 2'b01;
			14'b00101011110101: M1r = 2'b00;
			14'b01101011110101: M1r = 2'b01;
			14'b10101011110101: M1r = 2'b01;
			14'b11101011110101: M1r = 2'b01;
			14'b00111011110101: M1r = 2'b00;
			14'b01111011110101: M1r = 2'b00;
			14'b10111011110101: M1r = 2'b00;
			14'b11111011110101: M1r = 2'b00;
			14'b00001111110101: M1r = 2'b10;
			14'b01001111110101: M1r = 2'b10;
			14'b10001111110101: M1r = 2'b10;
			14'b11001111110101: M1r = 2'b11;
			14'b00011111110101: M1r = 2'b10;
			14'b01011111110101: M1r = 2'b10;
			14'b10011111110101: M1r = 2'b10;
			14'b11011111110101: M1r = 2'b10;
			14'b00101111110101: M1r = 2'b01;
			14'b01101111110101: M1r = 2'b01;
			14'b10101111110101: M1r = 2'b01;
			14'b11101111110101: M1r = 2'b10;
			14'b00111111110101: M1r = 2'b01;
			14'b01111111110101: M1r = 2'b01;
			14'b10111111110101: M1r = 2'b01;
			14'b11111111110101: M1r = 2'b01;
			14'b00000000001001: M1r = 2'b00;
			14'b01000000001001: M1r = 2'b00;
			14'b10000000001001: M1r = 2'b00;
			14'b11000000001001: M1r = 2'b00;
			14'b00010000001001: M1r = 2'b00;
			14'b01010000001001: M1r = 2'b00;
			14'b10010000001001: M1r = 2'b00;
			14'b11010000001001: M1r = 2'b00;
			14'b00100000001001: M1r = 2'b00;
			14'b01100000001001: M1r = 2'b00;
			14'b10100000001001: M1r = 2'b00;
			14'b11100000001001: M1r = 2'b00;
			14'b00110000001001: M1r = 2'b00;
			14'b01110000001001: M1r = 2'b00;
			14'b10110000001001: M1r = 2'b00;
			14'b11110000001001: M1r = 2'b00;
			14'b00000100001001: M1r = 2'b00;
			14'b01000100001001: M1r = 2'b00;
			14'b10000100001001: M1r = 2'b00;
			14'b11000100001001: M1r = 2'b00;
			14'b00010100001001: M1r = 2'b00;
			14'b01010100001001: M1r = 2'b00;
			14'b10010100001001: M1r = 2'b00;
			14'b11010100001001: M1r = 2'b00;
			14'b00100100001001: M1r = 2'b00;
			14'b01100100001001: M1r = 2'b00;
			14'b10100100001001: M1r = 2'b00;
			14'b11100100001001: M1r = 2'b00;
			14'b00110100001001: M1r = 2'b00;
			14'b01110100001001: M1r = 2'b00;
			14'b10110100001001: M1r = 2'b00;
			14'b11110100001001: M1r = 2'b00;
			14'b00001000001001: M1r = 2'b00;
			14'b01001000001001: M1r = 2'b00;
			14'b10001000001001: M1r = 2'b00;
			14'b11001000001001: M1r = 2'b01;
			14'b00011000001001: M1r = 2'b00;
			14'b01011000001001: M1r = 2'b00;
			14'b10011000001001: M1r = 2'b00;
			14'b11011000001001: M1r = 2'b00;
			14'b00101000001001: M1r = 2'b00;
			14'b01101000001001: M1r = 2'b00;
			14'b10101000001001: M1r = 2'b00;
			14'b11101000001001: M1r = 2'b00;
			14'b00111000001001: M1r = 2'b00;
			14'b01111000001001: M1r = 2'b00;
			14'b10111000001001: M1r = 2'b00;
			14'b11111000001001: M1r = 2'b00;
			14'b00001100001001: M1r = 2'b01;
			14'b01001100001001: M1r = 2'b01;
			14'b10001100001001: M1r = 2'b01;
			14'b11001100001001: M1r = 2'b01;
			14'b00011100001001: M1r = 2'b00;
			14'b01011100001001: M1r = 2'b00;
			14'b10011100001001: M1r = 2'b01;
			14'b11011100001001: M1r = 2'b01;
			14'b00101100001001: M1r = 2'b00;
			14'b01101100001001: M1r = 2'b00;
			14'b10101100001001: M1r = 2'b00;
			14'b11101100001001: M1r = 2'b00;
			14'b00111100001001: M1r = 2'b00;
			14'b01111100001001: M1r = 2'b00;
			14'b10111100001001: M1r = 2'b00;
			14'b11111100001001: M1r = 2'b00;
			14'b00000001001001: M1r = 2'b00;
			14'b01000001001001: M1r = 2'b00;
			14'b10000001001001: M1r = 2'b00;
			14'b11000001001001: M1r = 2'b00;
			14'b00010001001001: M1r = 2'b00;
			14'b01010001001001: M1r = 2'b00;
			14'b10010001001001: M1r = 2'b00;
			14'b11010001001001: M1r = 2'b00;
			14'b00100001001001: M1r = 2'b00;
			14'b01100001001001: M1r = 2'b00;
			14'b10100001001001: M1r = 2'b00;
			14'b11100001001001: M1r = 2'b00;
			14'b00110001001001: M1r = 2'b00;
			14'b01110001001001: M1r = 2'b00;
			14'b10110001001001: M1r = 2'b00;
			14'b11110001001001: M1r = 2'b00;
			14'b00000101001001: M1r = 2'b00;
			14'b01000101001001: M1r = 2'b00;
			14'b10000101001001: M1r = 2'b00;
			14'b11000101001001: M1r = 2'b00;
			14'b00010101001001: M1r = 2'b00;
			14'b01010101001001: M1r = 2'b00;
			14'b10010101001001: M1r = 2'b00;
			14'b11010101001001: M1r = 2'b00;
			14'b00100101001001: M1r = 2'b00;
			14'b01100101001001: M1r = 2'b00;
			14'b10100101001001: M1r = 2'b00;
			14'b11100101001001: M1r = 2'b00;
			14'b00110101001001: M1r = 2'b00;
			14'b01110101001001: M1r = 2'b00;
			14'b10110101001001: M1r = 2'b00;
			14'b11110101001001: M1r = 2'b00;
			14'b00001001001001: M1r = 2'b00;
			14'b01001001001001: M1r = 2'b00;
			14'b10001001001001: M1r = 2'b00;
			14'b11001001001001: M1r = 2'b00;
			14'b00011001001001: M1r = 2'b00;
			14'b01011001001001: M1r = 2'b00;
			14'b10011001001001: M1r = 2'b00;
			14'b11011001001001: M1r = 2'b00;
			14'b00101001001001: M1r = 2'b00;
			14'b01101001001001: M1r = 2'b00;
			14'b10101001001001: M1r = 2'b00;
			14'b11101001001001: M1r = 2'b00;
			14'b00111001001001: M1r = 2'b00;
			14'b01111001001001: M1r = 2'b00;
			14'b10111001001001: M1r = 2'b00;
			14'b11111001001001: M1r = 2'b00;
			14'b00001101001001: M1r = 2'b01;
			14'b01001101001001: M1r = 2'b01;
			14'b10001101001001: M1r = 2'b01;
			14'b11001101001001: M1r = 2'b01;
			14'b00011101001001: M1r = 2'b00;
			14'b01011101001001: M1r = 2'b00;
			14'b10011101001001: M1r = 2'b00;
			14'b11011101001001: M1r = 2'b01;
			14'b00101101001001: M1r = 2'b00;
			14'b01101101001001: M1r = 2'b00;
			14'b10101101001001: M1r = 2'b00;
			14'b11101101001001: M1r = 2'b00;
			14'b00111101001001: M1r = 2'b00;
			14'b01111101001001: M1r = 2'b00;
			14'b10111101001001: M1r = 2'b00;
			14'b11111101001001: M1r = 2'b00;
			14'b00000010001001: M1r = 2'b00;
			14'b01000010001001: M1r = 2'b00;
			14'b10000010001001: M1r = 2'b00;
			14'b11000010001001: M1r = 2'b00;
			14'b00010010001001: M1r = 2'b00;
			14'b01010010001001: M1r = 2'b00;
			14'b10010010001001: M1r = 2'b00;
			14'b11010010001001: M1r = 2'b00;
			14'b00100010001001: M1r = 2'b00;
			14'b01100010001001: M1r = 2'b00;
			14'b10100010001001: M1r = 2'b00;
			14'b11100010001001: M1r = 2'b00;
			14'b00110010001001: M1r = 2'b00;
			14'b01110010001001: M1r = 2'b00;
			14'b10110010001001: M1r = 2'b00;
			14'b11110010001001: M1r = 2'b00;
			14'b00000110001001: M1r = 2'b00;
			14'b01000110001001: M1r = 2'b00;
			14'b10000110001001: M1r = 2'b00;
			14'b11000110001001: M1r = 2'b00;
			14'b00010110001001: M1r = 2'b00;
			14'b01010110001001: M1r = 2'b00;
			14'b10010110001001: M1r = 2'b00;
			14'b11010110001001: M1r = 2'b00;
			14'b00100110001001: M1r = 2'b00;
			14'b01100110001001: M1r = 2'b00;
			14'b10100110001001: M1r = 2'b00;
			14'b11100110001001: M1r = 2'b00;
			14'b00110110001001: M1r = 2'b00;
			14'b01110110001001: M1r = 2'b00;
			14'b10110110001001: M1r = 2'b00;
			14'b11110110001001: M1r = 2'b00;
			14'b00001010001001: M1r = 2'b00;
			14'b01001010001001: M1r = 2'b00;
			14'b10001010001001: M1r = 2'b00;
			14'b11001010001001: M1r = 2'b00;
			14'b00011010001001: M1r = 2'b00;
			14'b01011010001001: M1r = 2'b00;
			14'b10011010001001: M1r = 2'b00;
			14'b11011010001001: M1r = 2'b00;
			14'b00101010001001: M1r = 2'b00;
			14'b01101010001001: M1r = 2'b00;
			14'b10101010001001: M1r = 2'b00;
			14'b11101010001001: M1r = 2'b00;
			14'b00111010001001: M1r = 2'b00;
			14'b01111010001001: M1r = 2'b00;
			14'b10111010001001: M1r = 2'b00;
			14'b11111010001001: M1r = 2'b00;
			14'b00001110001001: M1r = 2'b00;
			14'b01001110001001: M1r = 2'b00;
			14'b10001110001001: M1r = 2'b01;
			14'b11001110001001: M1r = 2'b01;
			14'b00011110001001: M1r = 2'b00;
			14'b01011110001001: M1r = 2'b00;
			14'b10011110001001: M1r = 2'b00;
			14'b11011110001001: M1r = 2'b00;
			14'b00101110001001: M1r = 2'b00;
			14'b01101110001001: M1r = 2'b00;
			14'b10101110001001: M1r = 2'b00;
			14'b11101110001001: M1r = 2'b00;
			14'b00111110001001: M1r = 2'b00;
			14'b01111110001001: M1r = 2'b00;
			14'b10111110001001: M1r = 2'b00;
			14'b11111110001001: M1r = 2'b00;
			14'b00000011001001: M1r = 2'b00;
			14'b01000011001001: M1r = 2'b00;
			14'b10000011001001: M1r = 2'b00;
			14'b11000011001001: M1r = 2'b00;
			14'b00010011001001: M1r = 2'b00;
			14'b01010011001001: M1r = 2'b00;
			14'b10010011001001: M1r = 2'b00;
			14'b11010011001001: M1r = 2'b00;
			14'b00100011001001: M1r = 2'b00;
			14'b01100011001001: M1r = 2'b00;
			14'b10100011001001: M1r = 2'b00;
			14'b11100011001001: M1r = 2'b00;
			14'b00110011001001: M1r = 2'b00;
			14'b01110011001001: M1r = 2'b00;
			14'b10110011001001: M1r = 2'b00;
			14'b11110011001001: M1r = 2'b00;
			14'b00000111001001: M1r = 2'b00;
			14'b01000111001001: M1r = 2'b00;
			14'b10000111001001: M1r = 2'b00;
			14'b11000111001001: M1r = 2'b00;
			14'b00010111001001: M1r = 2'b00;
			14'b01010111001001: M1r = 2'b00;
			14'b10010111001001: M1r = 2'b00;
			14'b11010111001001: M1r = 2'b00;
			14'b00100111001001: M1r = 2'b00;
			14'b01100111001001: M1r = 2'b00;
			14'b10100111001001: M1r = 2'b00;
			14'b11100111001001: M1r = 2'b00;
			14'b00110111001001: M1r = 2'b00;
			14'b01110111001001: M1r = 2'b00;
			14'b10110111001001: M1r = 2'b00;
			14'b11110111001001: M1r = 2'b00;
			14'b00001011001001: M1r = 2'b00;
			14'b01001011001001: M1r = 2'b00;
			14'b10001011001001: M1r = 2'b00;
			14'b11001011001001: M1r = 2'b00;
			14'b00011011001001: M1r = 2'b00;
			14'b01011011001001: M1r = 2'b00;
			14'b10011011001001: M1r = 2'b00;
			14'b11011011001001: M1r = 2'b00;
			14'b00101011001001: M1r = 2'b00;
			14'b01101011001001: M1r = 2'b00;
			14'b10101011001001: M1r = 2'b00;
			14'b11101011001001: M1r = 2'b00;
			14'b00111011001001: M1r = 2'b00;
			14'b01111011001001: M1r = 2'b00;
			14'b10111011001001: M1r = 2'b00;
			14'b11111011001001: M1r = 2'b00;
			14'b00001111001001: M1r = 2'b00;
			14'b01001111001001: M1r = 2'b00;
			14'b10001111001001: M1r = 2'b00;
			14'b11001111001001: M1r = 2'b00;
			14'b00011111001001: M1r = 2'b00;
			14'b01011111001001: M1r = 2'b00;
			14'b10011111001001: M1r = 2'b00;
			14'b11011111001001: M1r = 2'b00;
			14'b00101111001001: M1r = 2'b00;
			14'b01101111001001: M1r = 2'b00;
			14'b10101111001001: M1r = 2'b00;
			14'b11101111001001: M1r = 2'b00;
			14'b00111111001001: M1r = 2'b00;
			14'b01111111001001: M1r = 2'b00;
			14'b10111111001001: M1r = 2'b00;
			14'b11111111001001: M1r = 2'b00;
			14'b00000000011001: M1r = 2'b00;
			14'b01000000011001: M1r = 2'b00;
			14'b10000000011001: M1r = 2'b00;
			14'b11000000011001: M1r = 2'b00;
			14'b00010000011001: M1r = 2'b00;
			14'b01010000011001: M1r = 2'b00;
			14'b10010000011001: M1r = 2'b00;
			14'b11010000011001: M1r = 2'b00;
			14'b00100000011001: M1r = 2'b00;
			14'b01100000011001: M1r = 2'b00;
			14'b10100000011001: M1r = 2'b00;
			14'b11100000011001: M1r = 2'b00;
			14'b00110000011001: M1r = 2'b00;
			14'b01110000011001: M1r = 2'b00;
			14'b10110000011001: M1r = 2'b00;
			14'b11110000011001: M1r = 2'b00;
			14'b00000100011001: M1r = 2'b00;
			14'b01000100011001: M1r = 2'b00;
			14'b10000100011001: M1r = 2'b00;
			14'b11000100011001: M1r = 2'b00;
			14'b00010100011001: M1r = 2'b00;
			14'b01010100011001: M1r = 2'b00;
			14'b10010100011001: M1r = 2'b00;
			14'b11010100011001: M1r = 2'b00;
			14'b00100100011001: M1r = 2'b00;
			14'b01100100011001: M1r = 2'b00;
			14'b10100100011001: M1r = 2'b00;
			14'b11100100011001: M1r = 2'b00;
			14'b00110100011001: M1r = 2'b00;
			14'b01110100011001: M1r = 2'b00;
			14'b10110100011001: M1r = 2'b00;
			14'b11110100011001: M1r = 2'b00;
			14'b00001000011001: M1r = 2'b00;
			14'b01001000011001: M1r = 2'b01;
			14'b10001000011001: M1r = 2'b01;
			14'b11001000011001: M1r = 2'b01;
			14'b00011000011001: M1r = 2'b00;
			14'b01011000011001: M1r = 2'b00;
			14'b10011000011001: M1r = 2'b00;
			14'b11011000011001: M1r = 2'b00;
			14'b00101000011001: M1r = 2'b00;
			14'b01101000011001: M1r = 2'b00;
			14'b10101000011001: M1r = 2'b00;
			14'b11101000011001: M1r = 2'b00;
			14'b00111000011001: M1r = 2'b00;
			14'b01111000011001: M1r = 2'b00;
			14'b10111000011001: M1r = 2'b00;
			14'b11111000011001: M1r = 2'b00;
			14'b00001100011001: M1r = 2'b01;
			14'b01001100011001: M1r = 2'b01;
			14'b10001100011001: M1r = 2'b10;
			14'b11001100011001: M1r = 2'b10;
			14'b00011100011001: M1r = 2'b01;
			14'b01011100011001: M1r = 2'b01;
			14'b10011100011001: M1r = 2'b01;
			14'b11011100011001: M1r = 2'b01;
			14'b00101100011001: M1r = 2'b00;
			14'b01101100011001: M1r = 2'b00;
			14'b10101100011001: M1r = 2'b01;
			14'b11101100011001: M1r = 2'b01;
			14'b00111100011001: M1r = 2'b00;
			14'b01111100011001: M1r = 2'b00;
			14'b10111100011001: M1r = 2'b00;
			14'b11111100011001: M1r = 2'b00;
			14'b00000001011001: M1r = 2'b00;
			14'b01000001011001: M1r = 2'b00;
			14'b10000001011001: M1r = 2'b00;
			14'b11000001011001: M1r = 2'b00;
			14'b00010001011001: M1r = 2'b00;
			14'b01010001011001: M1r = 2'b00;
			14'b10010001011001: M1r = 2'b00;
			14'b11010001011001: M1r = 2'b00;
			14'b00100001011001: M1r = 2'b00;
			14'b01100001011001: M1r = 2'b00;
			14'b10100001011001: M1r = 2'b00;
			14'b11100001011001: M1r = 2'b00;
			14'b00110001011001: M1r = 2'b00;
			14'b01110001011001: M1r = 2'b00;
			14'b10110001011001: M1r = 2'b00;
			14'b11110001011001: M1r = 2'b00;
			14'b00000101011001: M1r = 2'b00;
			14'b01000101011001: M1r = 2'b00;
			14'b10000101011001: M1r = 2'b00;
			14'b11000101011001: M1r = 2'b00;
			14'b00010101011001: M1r = 2'b00;
			14'b01010101011001: M1r = 2'b00;
			14'b10010101011001: M1r = 2'b00;
			14'b11010101011001: M1r = 2'b00;
			14'b00100101011001: M1r = 2'b00;
			14'b01100101011001: M1r = 2'b00;
			14'b10100101011001: M1r = 2'b00;
			14'b11100101011001: M1r = 2'b00;
			14'b00110101011001: M1r = 2'b00;
			14'b01110101011001: M1r = 2'b00;
			14'b10110101011001: M1r = 2'b00;
			14'b11110101011001: M1r = 2'b00;
			14'b00001001011001: M1r = 2'b00;
			14'b01001001011001: M1r = 2'b00;
			14'b10001001011001: M1r = 2'b01;
			14'b11001001011001: M1r = 2'b01;
			14'b00011001011001: M1r = 2'b00;
			14'b01011001011001: M1r = 2'b00;
			14'b10011001011001: M1r = 2'b00;
			14'b11011001011001: M1r = 2'b00;
			14'b00101001011001: M1r = 2'b00;
			14'b01101001011001: M1r = 2'b00;
			14'b10101001011001: M1r = 2'b00;
			14'b11101001011001: M1r = 2'b00;
			14'b00111001011001: M1r = 2'b00;
			14'b01111001011001: M1r = 2'b00;
			14'b10111001011001: M1r = 2'b00;
			14'b11111001011001: M1r = 2'b00;
			14'b00001101011001: M1r = 2'b01;
			14'b01001101011001: M1r = 2'b01;
			14'b10001101011001: M1r = 2'b01;
			14'b11001101011001: M1r = 2'b01;
			14'b00011101011001: M1r = 2'b00;
			14'b01011101011001: M1r = 2'b01;
			14'b10011101011001: M1r = 2'b01;
			14'b11011101011001: M1r = 2'b01;
			14'b00101101011001: M1r = 2'b00;
			14'b01101101011001: M1r = 2'b00;
			14'b10101101011001: M1r = 2'b00;
			14'b11101101011001: M1r = 2'b00;
			14'b00111101011001: M1r = 2'b00;
			14'b01111101011001: M1r = 2'b00;
			14'b10111101011001: M1r = 2'b00;
			14'b11111101011001: M1r = 2'b00;
			14'b00000010011001: M1r = 2'b00;
			14'b01000010011001: M1r = 2'b00;
			14'b10000010011001: M1r = 2'b00;
			14'b11000010011001: M1r = 2'b00;
			14'b00010010011001: M1r = 2'b00;
			14'b01010010011001: M1r = 2'b00;
			14'b10010010011001: M1r = 2'b00;
			14'b11010010011001: M1r = 2'b00;
			14'b00100010011001: M1r = 2'b00;
			14'b01100010011001: M1r = 2'b00;
			14'b10100010011001: M1r = 2'b00;
			14'b11100010011001: M1r = 2'b00;
			14'b00110010011001: M1r = 2'b00;
			14'b01110010011001: M1r = 2'b00;
			14'b10110010011001: M1r = 2'b00;
			14'b11110010011001: M1r = 2'b00;
			14'b00000110011001: M1r = 2'b00;
			14'b01000110011001: M1r = 2'b00;
			14'b10000110011001: M1r = 2'b00;
			14'b11000110011001: M1r = 2'b00;
			14'b00010110011001: M1r = 2'b00;
			14'b01010110011001: M1r = 2'b00;
			14'b10010110011001: M1r = 2'b00;
			14'b11010110011001: M1r = 2'b00;
			14'b00100110011001: M1r = 2'b00;
			14'b01100110011001: M1r = 2'b00;
			14'b10100110011001: M1r = 2'b00;
			14'b11100110011001: M1r = 2'b00;
			14'b00110110011001: M1r = 2'b00;
			14'b01110110011001: M1r = 2'b00;
			14'b10110110011001: M1r = 2'b00;
			14'b11110110011001: M1r = 2'b00;
			14'b00001010011001: M1r = 2'b00;
			14'b01001010011001: M1r = 2'b00;
			14'b10001010011001: M1r = 2'b00;
			14'b11001010011001: M1r = 2'b00;
			14'b00011010011001: M1r = 2'b00;
			14'b01011010011001: M1r = 2'b00;
			14'b10011010011001: M1r = 2'b00;
			14'b11011010011001: M1r = 2'b00;
			14'b00101010011001: M1r = 2'b00;
			14'b01101010011001: M1r = 2'b00;
			14'b10101010011001: M1r = 2'b00;
			14'b11101010011001: M1r = 2'b00;
			14'b00111010011001: M1r = 2'b00;
			14'b01111010011001: M1r = 2'b00;
			14'b10111010011001: M1r = 2'b00;
			14'b11111010011001: M1r = 2'b00;
			14'b00001110011001: M1r = 2'b01;
			14'b01001110011001: M1r = 2'b01;
			14'b10001110011001: M1r = 2'b01;
			14'b11001110011001: M1r = 2'b01;
			14'b00011110011001: M1r = 2'b00;
			14'b01011110011001: M1r = 2'b00;
			14'b10011110011001: M1r = 2'b01;
			14'b11011110011001: M1r = 2'b01;
			14'b00101110011001: M1r = 2'b00;
			14'b01101110011001: M1r = 2'b00;
			14'b10101110011001: M1r = 2'b00;
			14'b11101110011001: M1r = 2'b00;
			14'b00111110011001: M1r = 2'b00;
			14'b01111110011001: M1r = 2'b00;
			14'b10111110011001: M1r = 2'b00;
			14'b11111110011001: M1r = 2'b00;
			14'b00000011011001: M1r = 2'b00;
			14'b01000011011001: M1r = 2'b00;
			14'b10000011011001: M1r = 2'b00;
			14'b11000011011001: M1r = 2'b00;
			14'b00010011011001: M1r = 2'b00;
			14'b01010011011001: M1r = 2'b00;
			14'b10010011011001: M1r = 2'b00;
			14'b11010011011001: M1r = 2'b00;
			14'b00100011011001: M1r = 2'b00;
			14'b01100011011001: M1r = 2'b00;
			14'b10100011011001: M1r = 2'b00;
			14'b11100011011001: M1r = 2'b00;
			14'b00110011011001: M1r = 2'b00;
			14'b01110011011001: M1r = 2'b00;
			14'b10110011011001: M1r = 2'b00;
			14'b11110011011001: M1r = 2'b00;
			14'b00000111011001: M1r = 2'b00;
			14'b01000111011001: M1r = 2'b00;
			14'b10000111011001: M1r = 2'b00;
			14'b11000111011001: M1r = 2'b00;
			14'b00010111011001: M1r = 2'b00;
			14'b01010111011001: M1r = 2'b00;
			14'b10010111011001: M1r = 2'b00;
			14'b11010111011001: M1r = 2'b00;
			14'b00100111011001: M1r = 2'b00;
			14'b01100111011001: M1r = 2'b00;
			14'b10100111011001: M1r = 2'b00;
			14'b11100111011001: M1r = 2'b00;
			14'b00110111011001: M1r = 2'b00;
			14'b01110111011001: M1r = 2'b00;
			14'b10110111011001: M1r = 2'b00;
			14'b11110111011001: M1r = 2'b00;
			14'b00001011011001: M1r = 2'b00;
			14'b01001011011001: M1r = 2'b00;
			14'b10001011011001: M1r = 2'b00;
			14'b11001011011001: M1r = 2'b00;
			14'b00011011011001: M1r = 2'b00;
			14'b01011011011001: M1r = 2'b00;
			14'b10011011011001: M1r = 2'b00;
			14'b11011011011001: M1r = 2'b00;
			14'b00101011011001: M1r = 2'b00;
			14'b01101011011001: M1r = 2'b00;
			14'b10101011011001: M1r = 2'b00;
			14'b11101011011001: M1r = 2'b00;
			14'b00111011011001: M1r = 2'b00;
			14'b01111011011001: M1r = 2'b00;
			14'b10111011011001: M1r = 2'b00;
			14'b11111011011001: M1r = 2'b00;
			14'b00001111011001: M1r = 2'b00;
			14'b01001111011001: M1r = 2'b01;
			14'b10001111011001: M1r = 2'b01;
			14'b11001111011001: M1r = 2'b01;
			14'b00011111011001: M1r = 2'b00;
			14'b01011111011001: M1r = 2'b00;
			14'b10011111011001: M1r = 2'b00;
			14'b11011111011001: M1r = 2'b00;
			14'b00101111011001: M1r = 2'b00;
			14'b01101111011001: M1r = 2'b00;
			14'b10101111011001: M1r = 2'b00;
			14'b11101111011001: M1r = 2'b00;
			14'b00111111011001: M1r = 2'b00;
			14'b01111111011001: M1r = 2'b00;
			14'b10111111011001: M1r = 2'b00;
			14'b11111111011001: M1r = 2'b00;
			14'b00000000101001: M1r = 2'b00;
			14'b01000000101001: M1r = 2'b00;
			14'b10000000101001: M1r = 2'b00;
			14'b11000000101001: M1r = 2'b00;
			14'b00010000101001: M1r = 2'b00;
			14'b01010000101001: M1r = 2'b00;
			14'b10010000101001: M1r = 2'b00;
			14'b11010000101001: M1r = 2'b00;
			14'b00100000101001: M1r = 2'b00;
			14'b01100000101001: M1r = 2'b00;
			14'b10100000101001: M1r = 2'b00;
			14'b11100000101001: M1r = 2'b00;
			14'b00110000101001: M1r = 2'b00;
			14'b01110000101001: M1r = 2'b00;
			14'b10110000101001: M1r = 2'b00;
			14'b11110000101001: M1r = 2'b00;
			14'b00000100101001: M1r = 2'b00;
			14'b01000100101001: M1r = 2'b00;
			14'b10000100101001: M1r = 2'b00;
			14'b11000100101001: M1r = 2'b01;
			14'b00010100101001: M1r = 2'b00;
			14'b01010100101001: M1r = 2'b00;
			14'b10010100101001: M1r = 2'b00;
			14'b11010100101001: M1r = 2'b00;
			14'b00100100101001: M1r = 2'b00;
			14'b01100100101001: M1r = 2'b00;
			14'b10100100101001: M1r = 2'b00;
			14'b11100100101001: M1r = 2'b00;
			14'b00110100101001: M1r = 2'b00;
			14'b01110100101001: M1r = 2'b00;
			14'b10110100101001: M1r = 2'b00;
			14'b11110100101001: M1r = 2'b00;
			14'b00001000101001: M1r = 2'b01;
			14'b01001000101001: M1r = 2'b01;
			14'b10001000101001: M1r = 2'b01;
			14'b11001000101001: M1r = 2'b01;
			14'b00011000101001: M1r = 2'b00;
			14'b01011000101001: M1r = 2'b01;
			14'b10011000101001: M1r = 2'b01;
			14'b11011000101001: M1r = 2'b01;
			14'b00101000101001: M1r = 2'b00;
			14'b01101000101001: M1r = 2'b00;
			14'b10101000101001: M1r = 2'b00;
			14'b11101000101001: M1r = 2'b00;
			14'b00111000101001: M1r = 2'b00;
			14'b01111000101001: M1r = 2'b00;
			14'b10111000101001: M1r = 2'b00;
			14'b11111000101001: M1r = 2'b00;
			14'b00001100101001: M1r = 2'b10;
			14'b01001100101001: M1r = 2'b10;
			14'b10001100101001: M1r = 2'b10;
			14'b11001100101001: M1r = 2'b10;
			14'b00011100101001: M1r = 2'b01;
			14'b01011100101001: M1r = 2'b01;
			14'b10011100101001: M1r = 2'b01;
			14'b11011100101001: M1r = 2'b10;
			14'b00101100101001: M1r = 2'b01;
			14'b01101100101001: M1r = 2'b01;
			14'b10101100101001: M1r = 2'b01;
			14'b11101100101001: M1r = 2'b01;
			14'b00111100101001: M1r = 2'b00;
			14'b01111100101001: M1r = 2'b00;
			14'b10111100101001: M1r = 2'b01;
			14'b11111100101001: M1r = 2'b01;
			14'b00000001101001: M1r = 2'b00;
			14'b01000001101001: M1r = 2'b00;
			14'b10000001101001: M1r = 2'b00;
			14'b11000001101001: M1r = 2'b00;
			14'b00010001101001: M1r = 2'b00;
			14'b01010001101001: M1r = 2'b00;
			14'b10010001101001: M1r = 2'b00;
			14'b11010001101001: M1r = 2'b00;
			14'b00100001101001: M1r = 2'b00;
			14'b01100001101001: M1r = 2'b00;
			14'b10100001101001: M1r = 2'b00;
			14'b11100001101001: M1r = 2'b00;
			14'b00110001101001: M1r = 2'b00;
			14'b01110001101001: M1r = 2'b00;
			14'b10110001101001: M1r = 2'b00;
			14'b11110001101001: M1r = 2'b00;
			14'b00000101101001: M1r = 2'b00;
			14'b01000101101001: M1r = 2'b00;
			14'b10000101101001: M1r = 2'b00;
			14'b11000101101001: M1r = 2'b00;
			14'b00010101101001: M1r = 2'b00;
			14'b01010101101001: M1r = 2'b00;
			14'b10010101101001: M1r = 2'b00;
			14'b11010101101001: M1r = 2'b00;
			14'b00100101101001: M1r = 2'b00;
			14'b01100101101001: M1r = 2'b00;
			14'b10100101101001: M1r = 2'b00;
			14'b11100101101001: M1r = 2'b00;
			14'b00110101101001: M1r = 2'b00;
			14'b01110101101001: M1r = 2'b00;
			14'b10110101101001: M1r = 2'b00;
			14'b11110101101001: M1r = 2'b00;
			14'b00001001101001: M1r = 2'b01;
			14'b01001001101001: M1r = 2'b01;
			14'b10001001101001: M1r = 2'b01;
			14'b11001001101001: M1r = 2'b01;
			14'b00011001101001: M1r = 2'b00;
			14'b01011001101001: M1r = 2'b00;
			14'b10011001101001: M1r = 2'b00;
			14'b11011001101001: M1r = 2'b01;
			14'b00101001101001: M1r = 2'b00;
			14'b01101001101001: M1r = 2'b00;
			14'b10101001101001: M1r = 2'b00;
			14'b11101001101001: M1r = 2'b00;
			14'b00111001101001: M1r = 2'b00;
			14'b01111001101001: M1r = 2'b00;
			14'b10111001101001: M1r = 2'b00;
			14'b11111001101001: M1r = 2'b00;
			14'b00001101101001: M1r = 2'b01;
			14'b01001101101001: M1r = 2'b10;
			14'b10001101101001: M1r = 2'b10;
			14'b11001101101001: M1r = 2'b10;
			14'b00011101101001: M1r = 2'b01;
			14'b01011101101001: M1r = 2'b01;
			14'b10011101101001: M1r = 2'b01;
			14'b11011101101001: M1r = 2'b01;
			14'b00101101101001: M1r = 2'b00;
			14'b01101101101001: M1r = 2'b01;
			14'b10101101101001: M1r = 2'b01;
			14'b11101101101001: M1r = 2'b01;
			14'b00111101101001: M1r = 2'b00;
			14'b01111101101001: M1r = 2'b00;
			14'b10111101101001: M1r = 2'b00;
			14'b11111101101001: M1r = 2'b00;
			14'b00000010101001: M1r = 2'b00;
			14'b01000010101001: M1r = 2'b00;
			14'b10000010101001: M1r = 2'b00;
			14'b11000010101001: M1r = 2'b00;
			14'b00010010101001: M1r = 2'b00;
			14'b01010010101001: M1r = 2'b00;
			14'b10010010101001: M1r = 2'b00;
			14'b11010010101001: M1r = 2'b00;
			14'b00100010101001: M1r = 2'b00;
			14'b01100010101001: M1r = 2'b00;
			14'b10100010101001: M1r = 2'b00;
			14'b11100010101001: M1r = 2'b00;
			14'b00110010101001: M1r = 2'b00;
			14'b01110010101001: M1r = 2'b00;
			14'b10110010101001: M1r = 2'b00;
			14'b11110010101001: M1r = 2'b00;
			14'b00000110101001: M1r = 2'b00;
			14'b01000110101001: M1r = 2'b00;
			14'b10000110101001: M1r = 2'b00;
			14'b11000110101001: M1r = 2'b00;
			14'b00010110101001: M1r = 2'b00;
			14'b01010110101001: M1r = 2'b00;
			14'b10010110101001: M1r = 2'b00;
			14'b11010110101001: M1r = 2'b00;
			14'b00100110101001: M1r = 2'b00;
			14'b01100110101001: M1r = 2'b00;
			14'b10100110101001: M1r = 2'b00;
			14'b11100110101001: M1r = 2'b00;
			14'b00110110101001: M1r = 2'b00;
			14'b01110110101001: M1r = 2'b00;
			14'b10110110101001: M1r = 2'b00;
			14'b11110110101001: M1r = 2'b00;
			14'b00001010101001: M1r = 2'b00;
			14'b01001010101001: M1r = 2'b01;
			14'b10001010101001: M1r = 2'b01;
			14'b11001010101001: M1r = 2'b01;
			14'b00011010101001: M1r = 2'b00;
			14'b01011010101001: M1r = 2'b00;
			14'b10011010101001: M1r = 2'b00;
			14'b11011010101001: M1r = 2'b00;
			14'b00101010101001: M1r = 2'b00;
			14'b01101010101001: M1r = 2'b00;
			14'b10101010101001: M1r = 2'b00;
			14'b11101010101001: M1r = 2'b00;
			14'b00111010101001: M1r = 2'b00;
			14'b01111010101001: M1r = 2'b00;
			14'b10111010101001: M1r = 2'b00;
			14'b11111010101001: M1r = 2'b00;
			14'b00001110101001: M1r = 2'b01;
			14'b01001110101001: M1r = 2'b01;
			14'b10001110101001: M1r = 2'b01;
			14'b11001110101001: M1r = 2'b10;
			14'b00011110101001: M1r = 2'b01;
			14'b01011110101001: M1r = 2'b01;
			14'b10011110101001: M1r = 2'b01;
			14'b11011110101001: M1r = 2'b01;
			14'b00101110101001: M1r = 2'b00;
			14'b01101110101001: M1r = 2'b00;
			14'b10101110101001: M1r = 2'b00;
			14'b11101110101001: M1r = 2'b01;
			14'b00111110101001: M1r = 2'b00;
			14'b01111110101001: M1r = 2'b00;
			14'b10111110101001: M1r = 2'b00;
			14'b11111110101001: M1r = 2'b00;
			14'b00000011101001: M1r = 2'b00;
			14'b01000011101001: M1r = 2'b00;
			14'b10000011101001: M1r = 2'b00;
			14'b11000011101001: M1r = 2'b00;
			14'b00010011101001: M1r = 2'b00;
			14'b01010011101001: M1r = 2'b00;
			14'b10010011101001: M1r = 2'b00;
			14'b11010011101001: M1r = 2'b00;
			14'b00100011101001: M1r = 2'b00;
			14'b01100011101001: M1r = 2'b00;
			14'b10100011101001: M1r = 2'b00;
			14'b11100011101001: M1r = 2'b00;
			14'b00110011101001: M1r = 2'b00;
			14'b01110011101001: M1r = 2'b00;
			14'b10110011101001: M1r = 2'b00;
			14'b11110011101001: M1r = 2'b00;
			14'b00000111101001: M1r = 2'b00;
			14'b01000111101001: M1r = 2'b00;
			14'b10000111101001: M1r = 2'b00;
			14'b11000111101001: M1r = 2'b00;
			14'b00010111101001: M1r = 2'b00;
			14'b01010111101001: M1r = 2'b00;
			14'b10010111101001: M1r = 2'b00;
			14'b11010111101001: M1r = 2'b00;
			14'b00100111101001: M1r = 2'b00;
			14'b01100111101001: M1r = 2'b00;
			14'b10100111101001: M1r = 2'b00;
			14'b11100111101001: M1r = 2'b00;
			14'b00110111101001: M1r = 2'b00;
			14'b01110111101001: M1r = 2'b00;
			14'b10110111101001: M1r = 2'b00;
			14'b11110111101001: M1r = 2'b00;
			14'b00001011101001: M1r = 2'b00;
			14'b01001011101001: M1r = 2'b00;
			14'b10001011101001: M1r = 2'b00;
			14'b11001011101001: M1r = 2'b01;
			14'b00011011101001: M1r = 2'b00;
			14'b01011011101001: M1r = 2'b00;
			14'b10011011101001: M1r = 2'b00;
			14'b11011011101001: M1r = 2'b00;
			14'b00101011101001: M1r = 2'b00;
			14'b01101011101001: M1r = 2'b00;
			14'b10101011101001: M1r = 2'b00;
			14'b11101011101001: M1r = 2'b00;
			14'b00111011101001: M1r = 2'b00;
			14'b01111011101001: M1r = 2'b00;
			14'b10111011101001: M1r = 2'b00;
			14'b11111011101001: M1r = 2'b00;
			14'b00001111101001: M1r = 2'b01;
			14'b01001111101001: M1r = 2'b01;
			14'b10001111101001: M1r = 2'b01;
			14'b11001111101001: M1r = 2'b01;
			14'b00011111101001: M1r = 2'b00;
			14'b01011111101001: M1r = 2'b01;
			14'b10011111101001: M1r = 2'b01;
			14'b11011111101001: M1r = 2'b01;
			14'b00101111101001: M1r = 2'b00;
			14'b01101111101001: M1r = 2'b00;
			14'b10101111101001: M1r = 2'b00;
			14'b11101111101001: M1r = 2'b00;
			14'b00111111101001: M1r = 2'b00;
			14'b01111111101001: M1r = 2'b00;
			14'b10111111101001: M1r = 2'b00;
			14'b11111111101001: M1r = 2'b00;
			14'b00000000111001: M1r = 2'b00;
			14'b01000000111001: M1r = 2'b00;
			14'b10000000111001: M1r = 2'b00;
			14'b11000000111001: M1r = 2'b00;
			14'b00010000111001: M1r = 2'b00;
			14'b01010000111001: M1r = 2'b00;
			14'b10010000111001: M1r = 2'b00;
			14'b11010000111001: M1r = 2'b00;
			14'b00100000111001: M1r = 2'b00;
			14'b01100000111001: M1r = 2'b00;
			14'b10100000111001: M1r = 2'b00;
			14'b11100000111001: M1r = 2'b00;
			14'b00110000111001: M1r = 2'b00;
			14'b01110000111001: M1r = 2'b00;
			14'b10110000111001: M1r = 2'b00;
			14'b11110000111001: M1r = 2'b00;
			14'b00000100111001: M1r = 2'b01;
			14'b01000100111001: M1r = 2'b01;
			14'b10000100111001: M1r = 2'b01;
			14'b11000100111001: M1r = 2'b01;
			14'b00010100111001: M1r = 2'b00;
			14'b01010100111001: M1r = 2'b00;
			14'b10010100111001: M1r = 2'b00;
			14'b11010100111001: M1r = 2'b01;
			14'b00100100111001: M1r = 2'b00;
			14'b01100100111001: M1r = 2'b00;
			14'b10100100111001: M1r = 2'b00;
			14'b11100100111001: M1r = 2'b00;
			14'b00110100111001: M1r = 2'b00;
			14'b01110100111001: M1r = 2'b00;
			14'b10110100111001: M1r = 2'b00;
			14'b11110100111001: M1r = 2'b00;
			14'b00001000111001: M1r = 2'b01;
			14'b01001000111001: M1r = 2'b01;
			14'b10001000111001: M1r = 2'b10;
			14'b11001000111001: M1r = 2'b10;
			14'b00011000111001: M1r = 2'b01;
			14'b01011000111001: M1r = 2'b01;
			14'b10011000111001: M1r = 2'b01;
			14'b11011000111001: M1r = 2'b01;
			14'b00101000111001: M1r = 2'b00;
			14'b01101000111001: M1r = 2'b01;
			14'b10101000111001: M1r = 2'b01;
			14'b11101000111001: M1r = 2'b01;
			14'b00111000111001: M1r = 2'b00;
			14'b01111000111001: M1r = 2'b00;
			14'b10111000111001: M1r = 2'b00;
			14'b11111000111001: M1r = 2'b00;
			14'b00001100111001: M1r = 2'b10;
			14'b01001100111001: M1r = 2'b10;
			14'b10001100111001: M1r = 2'b10;
			14'b11001100111001: M1r = 2'b11;
			14'b00011100111001: M1r = 2'b10;
			14'b01011100111001: M1r = 2'b10;
			14'b10011100111001: M1r = 2'b10;
			14'b11011100111001: M1r = 2'b10;
			14'b00101100111001: M1r = 2'b01;
			14'b01101100111001: M1r = 2'b01;
			14'b10101100111001: M1r = 2'b01;
			14'b11101100111001: M1r = 2'b10;
			14'b00111100111001: M1r = 2'b01;
			14'b01111100111001: M1r = 2'b01;
			14'b10111100111001: M1r = 2'b01;
			14'b11111100111001: M1r = 2'b01;
			14'b00000001111001: M1r = 2'b00;
			14'b01000001111001: M1r = 2'b00;
			14'b10000001111001: M1r = 2'b00;
			14'b11000001111001: M1r = 2'b00;
			14'b00010001111001: M1r = 2'b00;
			14'b01010001111001: M1r = 2'b00;
			14'b10010001111001: M1r = 2'b00;
			14'b11010001111001: M1r = 2'b00;
			14'b00100001111001: M1r = 2'b00;
			14'b01100001111001: M1r = 2'b00;
			14'b10100001111001: M1r = 2'b00;
			14'b11100001111001: M1r = 2'b00;
			14'b00110001111001: M1r = 2'b00;
			14'b01110001111001: M1r = 2'b00;
			14'b10110001111001: M1r = 2'b00;
			14'b11110001111001: M1r = 2'b00;
			14'b00000101111001: M1r = 2'b00;
			14'b01000101111001: M1r = 2'b00;
			14'b10000101111001: M1r = 2'b01;
			14'b11000101111001: M1r = 2'b01;
			14'b00010101111001: M1r = 2'b00;
			14'b01010101111001: M1r = 2'b00;
			14'b10010101111001: M1r = 2'b00;
			14'b11010101111001: M1r = 2'b00;
			14'b00100101111001: M1r = 2'b00;
			14'b01100101111001: M1r = 2'b00;
			14'b10100101111001: M1r = 2'b00;
			14'b11100101111001: M1r = 2'b00;
			14'b00110101111001: M1r = 2'b00;
			14'b01110101111001: M1r = 2'b00;
			14'b10110101111001: M1r = 2'b00;
			14'b11110101111001: M1r = 2'b00;
			14'b00001001111001: M1r = 2'b01;
			14'b01001001111001: M1r = 2'b01;
			14'b10001001111001: M1r = 2'b01;
			14'b11001001111001: M1r = 2'b10;
			14'b00011001111001: M1r = 2'b01;
			14'b01011001111001: M1r = 2'b01;
			14'b10011001111001: M1r = 2'b01;
			14'b11011001111001: M1r = 2'b01;
			14'b00101001111001: M1r = 2'b00;
			14'b01101001111001: M1r = 2'b00;
			14'b10101001111001: M1r = 2'b00;
			14'b11101001111001: M1r = 2'b01;
			14'b00111001111001: M1r = 2'b00;
			14'b01111001111001: M1r = 2'b00;
			14'b10111001111001: M1r = 2'b00;
			14'b11111001111001: M1r = 2'b00;
			14'b00001101111001: M1r = 2'b10;
			14'b01001101111001: M1r = 2'b10;
			14'b10001101111001: M1r = 2'b10;
			14'b11001101111001: M1r = 2'b10;
			14'b00011101111001: M1r = 2'b01;
			14'b01011101111001: M1r = 2'b01;
			14'b10011101111001: M1r = 2'b10;
			14'b11011101111001: M1r = 2'b10;
			14'b00101101111001: M1r = 2'b01;
			14'b01101101111001: M1r = 2'b01;
			14'b10101101111001: M1r = 2'b01;
			14'b11101101111001: M1r = 2'b01;
			14'b00111101111001: M1r = 2'b00;
			14'b01111101111001: M1r = 2'b01;
			14'b10111101111001: M1r = 2'b01;
			14'b11111101111001: M1r = 2'b01;
			14'b00000010111001: M1r = 2'b00;
			14'b01000010111001: M1r = 2'b00;
			14'b10000010111001: M1r = 2'b00;
			14'b11000010111001: M1r = 2'b00;
			14'b00010010111001: M1r = 2'b00;
			14'b01010010111001: M1r = 2'b00;
			14'b10010010111001: M1r = 2'b00;
			14'b11010010111001: M1r = 2'b00;
			14'b00100010111001: M1r = 2'b00;
			14'b01100010111001: M1r = 2'b00;
			14'b10100010111001: M1r = 2'b00;
			14'b11100010111001: M1r = 2'b00;
			14'b00110010111001: M1r = 2'b00;
			14'b01110010111001: M1r = 2'b00;
			14'b10110010111001: M1r = 2'b00;
			14'b11110010111001: M1r = 2'b00;
			14'b00000110111001: M1r = 2'b00;
			14'b01000110111001: M1r = 2'b00;
			14'b10000110111001: M1r = 2'b00;
			14'b11000110111001: M1r = 2'b01;
			14'b00010110111001: M1r = 2'b00;
			14'b01010110111001: M1r = 2'b00;
			14'b10010110111001: M1r = 2'b00;
			14'b11010110111001: M1r = 2'b00;
			14'b00100110111001: M1r = 2'b00;
			14'b01100110111001: M1r = 2'b00;
			14'b10100110111001: M1r = 2'b00;
			14'b11100110111001: M1r = 2'b00;
			14'b00110110111001: M1r = 2'b00;
			14'b01110110111001: M1r = 2'b00;
			14'b10110110111001: M1r = 2'b00;
			14'b11110110111001: M1r = 2'b00;
			14'b00001010111001: M1r = 2'b01;
			14'b01001010111001: M1r = 2'b01;
			14'b10001010111001: M1r = 2'b01;
			14'b11001010111001: M1r = 2'b01;
			14'b00011010111001: M1r = 2'b00;
			14'b01011010111001: M1r = 2'b00;
			14'b10011010111001: M1r = 2'b01;
			14'b11011010111001: M1r = 2'b01;
			14'b00101010111001: M1r = 2'b00;
			14'b01101010111001: M1r = 2'b00;
			14'b10101010111001: M1r = 2'b00;
			14'b11101010111001: M1r = 2'b00;
			14'b00111010111001: M1r = 2'b00;
			14'b01111010111001: M1r = 2'b00;
			14'b10111010111001: M1r = 2'b00;
			14'b11111010111001: M1r = 2'b00;
			14'b00001110111001: M1r = 2'b10;
			14'b01001110111001: M1r = 2'b10;
			14'b10001110111001: M1r = 2'b10;
			14'b11001110111001: M1r = 2'b10;
			14'b00011110111001: M1r = 2'b01;
			14'b01011110111001: M1r = 2'b01;
			14'b10011110111001: M1r = 2'b01;
			14'b11011110111001: M1r = 2'b10;
			14'b00101110111001: M1r = 2'b01;
			14'b01101110111001: M1r = 2'b01;
			14'b10101110111001: M1r = 2'b01;
			14'b11101110111001: M1r = 2'b01;
			14'b00111110111001: M1r = 2'b00;
			14'b01111110111001: M1r = 2'b00;
			14'b10111110111001: M1r = 2'b00;
			14'b11111110111001: M1r = 2'b01;
			14'b00000011111001: M1r = 2'b00;
			14'b01000011111001: M1r = 2'b00;
			14'b10000011111001: M1r = 2'b00;
			14'b11000011111001: M1r = 2'b00;
			14'b00010011111001: M1r = 2'b00;
			14'b01010011111001: M1r = 2'b00;
			14'b10010011111001: M1r = 2'b00;
			14'b11010011111001: M1r = 2'b00;
			14'b00100011111001: M1r = 2'b00;
			14'b01100011111001: M1r = 2'b00;
			14'b10100011111001: M1r = 2'b00;
			14'b11100011111001: M1r = 2'b00;
			14'b00110011111001: M1r = 2'b00;
			14'b01110011111001: M1r = 2'b00;
			14'b10110011111001: M1r = 2'b00;
			14'b11110011111001: M1r = 2'b00;
			14'b00000111111001: M1r = 2'b00;
			14'b01000111111001: M1r = 2'b00;
			14'b10000111111001: M1r = 2'b00;
			14'b11000111111001: M1r = 2'b00;
			14'b00010111111001: M1r = 2'b00;
			14'b01010111111001: M1r = 2'b00;
			14'b10010111111001: M1r = 2'b00;
			14'b11010111111001: M1r = 2'b00;
			14'b00100111111001: M1r = 2'b00;
			14'b01100111111001: M1r = 2'b00;
			14'b10100111111001: M1r = 2'b00;
			14'b11100111111001: M1r = 2'b00;
			14'b00110111111001: M1r = 2'b00;
			14'b01110111111001: M1r = 2'b00;
			14'b10110111111001: M1r = 2'b00;
			14'b11110111111001: M1r = 2'b00;
			14'b00001011111001: M1r = 2'b01;
			14'b01001011111001: M1r = 2'b01;
			14'b10001011111001: M1r = 2'b01;
			14'b11001011111001: M1r = 2'b01;
			14'b00011011111001: M1r = 2'b00;
			14'b01011011111001: M1r = 2'b00;
			14'b10011011111001: M1r = 2'b00;
			14'b11011011111001: M1r = 2'b01;
			14'b00101011111001: M1r = 2'b00;
			14'b01101011111001: M1r = 2'b00;
			14'b10101011111001: M1r = 2'b00;
			14'b11101011111001: M1r = 2'b00;
			14'b00111011111001: M1r = 2'b00;
			14'b01111011111001: M1r = 2'b00;
			14'b10111011111001: M1r = 2'b00;
			14'b11111011111001: M1r = 2'b00;
			14'b00001111111001: M1r = 2'b01;
			14'b01001111111001: M1r = 2'b01;
			14'b10001111111001: M1r = 2'b10;
			14'b11001111111001: M1r = 2'b10;
			14'b00011111111001: M1r = 2'b01;
			14'b01011111111001: M1r = 2'b01;
			14'b10011111111001: M1r = 2'b01;
			14'b11011111111001: M1r = 2'b01;
			14'b00101111111001: M1r = 2'b00;
			14'b01101111111001: M1r = 2'b00;
			14'b10101111111001: M1r = 2'b01;
			14'b11101111111001: M1r = 2'b01;
			14'b00111111111001: M1r = 2'b00;
			14'b01111111111001: M1r = 2'b00;
			14'b10111111111001: M1r = 2'b00;
			14'b11111111111001: M1r = 2'b00;
			14'b00000000001101: M1r = 2'b00;
			14'b01000000001101: M1r = 2'b00;
			14'b10000000001101: M1r = 2'b00;
			14'b11000000001101: M1r = 2'b00;
			14'b00010000001101: M1r = 2'b00;
			14'b01010000001101: M1r = 2'b00;
			14'b10010000001101: M1r = 2'b00;
			14'b11010000001101: M1r = 2'b00;
			14'b00100000001101: M1r = 2'b00;
			14'b01100000001101: M1r = 2'b00;
			14'b10100000001101: M1r = 2'b00;
			14'b11100000001101: M1r = 2'b00;
			14'b00110000001101: M1r = 2'b00;
			14'b01110000001101: M1r = 2'b00;
			14'b10110000001101: M1r = 2'b00;
			14'b11110000001101: M1r = 2'b00;
			14'b00000100001101: M1r = 2'b00;
			14'b01000100001101: M1r = 2'b00;
			14'b10000100001101: M1r = 2'b00;
			14'b11000100001101: M1r = 2'b00;
			14'b00010100001101: M1r = 2'b00;
			14'b01010100001101: M1r = 2'b00;
			14'b10010100001101: M1r = 2'b00;
			14'b11010100001101: M1r = 2'b00;
			14'b00100100001101: M1r = 2'b00;
			14'b01100100001101: M1r = 2'b00;
			14'b10100100001101: M1r = 2'b00;
			14'b11100100001101: M1r = 2'b00;
			14'b00110100001101: M1r = 2'b00;
			14'b01110100001101: M1r = 2'b00;
			14'b10110100001101: M1r = 2'b00;
			14'b11110100001101: M1r = 2'b00;
			14'b00001000001101: M1r = 2'b00;
			14'b01001000001101: M1r = 2'b00;
			14'b10001000001101: M1r = 2'b00;
			14'b11001000001101: M1r = 2'b00;
			14'b00011000001101: M1r = 2'b00;
			14'b01011000001101: M1r = 2'b00;
			14'b10011000001101: M1r = 2'b00;
			14'b11011000001101: M1r = 2'b00;
			14'b00101000001101: M1r = 2'b00;
			14'b01101000001101: M1r = 2'b00;
			14'b10101000001101: M1r = 2'b00;
			14'b11101000001101: M1r = 2'b00;
			14'b00111000001101: M1r = 2'b00;
			14'b01111000001101: M1r = 2'b00;
			14'b10111000001101: M1r = 2'b00;
			14'b11111000001101: M1r = 2'b00;
			14'b00001100001101: M1r = 2'b00;
			14'b01001100001101: M1r = 2'b00;
			14'b10001100001101: M1r = 2'b00;
			14'b11001100001101: M1r = 2'b00;
			14'b00011100001101: M1r = 2'b00;
			14'b01011100001101: M1r = 2'b00;
			14'b10011100001101: M1r = 2'b00;
			14'b11011100001101: M1r = 2'b00;
			14'b00101100001101: M1r = 2'b00;
			14'b01101100001101: M1r = 2'b00;
			14'b10101100001101: M1r = 2'b00;
			14'b11101100001101: M1r = 2'b00;
			14'b00111100001101: M1r = 2'b00;
			14'b01111100001101: M1r = 2'b00;
			14'b10111100001101: M1r = 2'b00;
			14'b11111100001101: M1r = 2'b00;
			14'b00000001001101: M1r = 2'b00;
			14'b01000001001101: M1r = 2'b00;
			14'b10000001001101: M1r = 2'b00;
			14'b11000001001101: M1r = 2'b00;
			14'b00010001001101: M1r = 2'b00;
			14'b01010001001101: M1r = 2'b00;
			14'b10010001001101: M1r = 2'b00;
			14'b11010001001101: M1r = 2'b00;
			14'b00100001001101: M1r = 2'b00;
			14'b01100001001101: M1r = 2'b00;
			14'b10100001001101: M1r = 2'b00;
			14'b11100001001101: M1r = 2'b00;
			14'b00110001001101: M1r = 2'b00;
			14'b01110001001101: M1r = 2'b00;
			14'b10110001001101: M1r = 2'b00;
			14'b11110001001101: M1r = 2'b00;
			14'b00000101001101: M1r = 2'b00;
			14'b01000101001101: M1r = 2'b00;
			14'b10000101001101: M1r = 2'b00;
			14'b11000101001101: M1r = 2'b00;
			14'b00010101001101: M1r = 2'b00;
			14'b01010101001101: M1r = 2'b00;
			14'b10010101001101: M1r = 2'b00;
			14'b11010101001101: M1r = 2'b00;
			14'b00100101001101: M1r = 2'b00;
			14'b01100101001101: M1r = 2'b00;
			14'b10100101001101: M1r = 2'b00;
			14'b11100101001101: M1r = 2'b00;
			14'b00110101001101: M1r = 2'b00;
			14'b01110101001101: M1r = 2'b00;
			14'b10110101001101: M1r = 2'b00;
			14'b11110101001101: M1r = 2'b00;
			14'b00001001001101: M1r = 2'b00;
			14'b01001001001101: M1r = 2'b00;
			14'b10001001001101: M1r = 2'b00;
			14'b11001001001101: M1r = 2'b00;
			14'b00011001001101: M1r = 2'b00;
			14'b01011001001101: M1r = 2'b00;
			14'b10011001001101: M1r = 2'b00;
			14'b11011001001101: M1r = 2'b00;
			14'b00101001001101: M1r = 2'b00;
			14'b01101001001101: M1r = 2'b00;
			14'b10101001001101: M1r = 2'b00;
			14'b11101001001101: M1r = 2'b00;
			14'b00111001001101: M1r = 2'b00;
			14'b01111001001101: M1r = 2'b00;
			14'b10111001001101: M1r = 2'b00;
			14'b11111001001101: M1r = 2'b00;
			14'b00001101001101: M1r = 2'b00;
			14'b01001101001101: M1r = 2'b00;
			14'b10001101001101: M1r = 2'b00;
			14'b11001101001101: M1r = 2'b00;
			14'b00011101001101: M1r = 2'b00;
			14'b01011101001101: M1r = 2'b00;
			14'b10011101001101: M1r = 2'b00;
			14'b11011101001101: M1r = 2'b00;
			14'b00101101001101: M1r = 2'b00;
			14'b01101101001101: M1r = 2'b00;
			14'b10101101001101: M1r = 2'b00;
			14'b11101101001101: M1r = 2'b00;
			14'b00111101001101: M1r = 2'b00;
			14'b01111101001101: M1r = 2'b00;
			14'b10111101001101: M1r = 2'b00;
			14'b11111101001101: M1r = 2'b00;
			14'b00000010001101: M1r = 2'b00;
			14'b01000010001101: M1r = 2'b00;
			14'b10000010001101: M1r = 2'b00;
			14'b11000010001101: M1r = 2'b00;
			14'b00010010001101: M1r = 2'b00;
			14'b01010010001101: M1r = 2'b00;
			14'b10010010001101: M1r = 2'b00;
			14'b11010010001101: M1r = 2'b00;
			14'b00100010001101: M1r = 2'b00;
			14'b01100010001101: M1r = 2'b00;
			14'b10100010001101: M1r = 2'b00;
			14'b11100010001101: M1r = 2'b00;
			14'b00110010001101: M1r = 2'b00;
			14'b01110010001101: M1r = 2'b00;
			14'b10110010001101: M1r = 2'b00;
			14'b11110010001101: M1r = 2'b00;
			14'b00000110001101: M1r = 2'b00;
			14'b01000110001101: M1r = 2'b00;
			14'b10000110001101: M1r = 2'b00;
			14'b11000110001101: M1r = 2'b00;
			14'b00010110001101: M1r = 2'b00;
			14'b01010110001101: M1r = 2'b00;
			14'b10010110001101: M1r = 2'b00;
			14'b11010110001101: M1r = 2'b00;
			14'b00100110001101: M1r = 2'b00;
			14'b01100110001101: M1r = 2'b00;
			14'b10100110001101: M1r = 2'b00;
			14'b11100110001101: M1r = 2'b00;
			14'b00110110001101: M1r = 2'b00;
			14'b01110110001101: M1r = 2'b00;
			14'b10110110001101: M1r = 2'b00;
			14'b11110110001101: M1r = 2'b00;
			14'b00001010001101: M1r = 2'b00;
			14'b01001010001101: M1r = 2'b00;
			14'b10001010001101: M1r = 2'b00;
			14'b11001010001101: M1r = 2'b00;
			14'b00011010001101: M1r = 2'b00;
			14'b01011010001101: M1r = 2'b00;
			14'b10011010001101: M1r = 2'b00;
			14'b11011010001101: M1r = 2'b00;
			14'b00101010001101: M1r = 2'b00;
			14'b01101010001101: M1r = 2'b00;
			14'b10101010001101: M1r = 2'b00;
			14'b11101010001101: M1r = 2'b00;
			14'b00111010001101: M1r = 2'b00;
			14'b01111010001101: M1r = 2'b00;
			14'b10111010001101: M1r = 2'b00;
			14'b11111010001101: M1r = 2'b00;
			14'b00001110001101: M1r = 2'b00;
			14'b01001110001101: M1r = 2'b00;
			14'b10001110001101: M1r = 2'b00;
			14'b11001110001101: M1r = 2'b00;
			14'b00011110001101: M1r = 2'b00;
			14'b01011110001101: M1r = 2'b00;
			14'b10011110001101: M1r = 2'b00;
			14'b11011110001101: M1r = 2'b00;
			14'b00101110001101: M1r = 2'b00;
			14'b01101110001101: M1r = 2'b00;
			14'b10101110001101: M1r = 2'b00;
			14'b11101110001101: M1r = 2'b00;
			14'b00111110001101: M1r = 2'b00;
			14'b01111110001101: M1r = 2'b00;
			14'b10111110001101: M1r = 2'b00;
			14'b11111110001101: M1r = 2'b00;
			14'b00000011001101: M1r = 2'b00;
			14'b01000011001101: M1r = 2'b00;
			14'b10000011001101: M1r = 2'b00;
			14'b11000011001101: M1r = 2'b00;
			14'b00010011001101: M1r = 2'b00;
			14'b01010011001101: M1r = 2'b00;
			14'b10010011001101: M1r = 2'b00;
			14'b11010011001101: M1r = 2'b00;
			14'b00100011001101: M1r = 2'b00;
			14'b01100011001101: M1r = 2'b00;
			14'b10100011001101: M1r = 2'b00;
			14'b11100011001101: M1r = 2'b00;
			14'b00110011001101: M1r = 2'b00;
			14'b01110011001101: M1r = 2'b00;
			14'b10110011001101: M1r = 2'b00;
			14'b11110011001101: M1r = 2'b00;
			14'b00000111001101: M1r = 2'b00;
			14'b01000111001101: M1r = 2'b00;
			14'b10000111001101: M1r = 2'b00;
			14'b11000111001101: M1r = 2'b00;
			14'b00010111001101: M1r = 2'b00;
			14'b01010111001101: M1r = 2'b00;
			14'b10010111001101: M1r = 2'b00;
			14'b11010111001101: M1r = 2'b00;
			14'b00100111001101: M1r = 2'b00;
			14'b01100111001101: M1r = 2'b00;
			14'b10100111001101: M1r = 2'b00;
			14'b11100111001101: M1r = 2'b00;
			14'b00110111001101: M1r = 2'b00;
			14'b01110111001101: M1r = 2'b00;
			14'b10110111001101: M1r = 2'b00;
			14'b11110111001101: M1r = 2'b00;
			14'b00001011001101: M1r = 2'b00;
			14'b01001011001101: M1r = 2'b00;
			14'b10001011001101: M1r = 2'b00;
			14'b11001011001101: M1r = 2'b00;
			14'b00011011001101: M1r = 2'b00;
			14'b01011011001101: M1r = 2'b00;
			14'b10011011001101: M1r = 2'b00;
			14'b11011011001101: M1r = 2'b00;
			14'b00101011001101: M1r = 2'b00;
			14'b01101011001101: M1r = 2'b00;
			14'b10101011001101: M1r = 2'b00;
			14'b11101011001101: M1r = 2'b00;
			14'b00111011001101: M1r = 2'b00;
			14'b01111011001101: M1r = 2'b00;
			14'b10111011001101: M1r = 2'b00;
			14'b11111011001101: M1r = 2'b00;
			14'b00001111001101: M1r = 2'b00;
			14'b01001111001101: M1r = 2'b00;
			14'b10001111001101: M1r = 2'b00;
			14'b11001111001101: M1r = 2'b00;
			14'b00011111001101: M1r = 2'b00;
			14'b01011111001101: M1r = 2'b00;
			14'b10011111001101: M1r = 2'b00;
			14'b11011111001101: M1r = 2'b00;
			14'b00101111001101: M1r = 2'b00;
			14'b01101111001101: M1r = 2'b00;
			14'b10101111001101: M1r = 2'b00;
			14'b11101111001101: M1r = 2'b00;
			14'b00111111001101: M1r = 2'b00;
			14'b01111111001101: M1r = 2'b00;
			14'b10111111001101: M1r = 2'b00;
			14'b11111111001101: M1r = 2'b00;
			14'b00000000011101: M1r = 2'b00;
			14'b01000000011101: M1r = 2'b00;
			14'b10000000011101: M1r = 2'b00;
			14'b11000000011101: M1r = 2'b00;
			14'b00010000011101: M1r = 2'b00;
			14'b01010000011101: M1r = 2'b00;
			14'b10010000011101: M1r = 2'b00;
			14'b11010000011101: M1r = 2'b00;
			14'b00100000011101: M1r = 2'b00;
			14'b01100000011101: M1r = 2'b00;
			14'b10100000011101: M1r = 2'b00;
			14'b11100000011101: M1r = 2'b00;
			14'b00110000011101: M1r = 2'b00;
			14'b01110000011101: M1r = 2'b00;
			14'b10110000011101: M1r = 2'b00;
			14'b11110000011101: M1r = 2'b00;
			14'b00000100011101: M1r = 2'b00;
			14'b01000100011101: M1r = 2'b00;
			14'b10000100011101: M1r = 2'b00;
			14'b11000100011101: M1r = 2'b00;
			14'b00010100011101: M1r = 2'b00;
			14'b01010100011101: M1r = 2'b00;
			14'b10010100011101: M1r = 2'b00;
			14'b11010100011101: M1r = 2'b00;
			14'b00100100011101: M1r = 2'b00;
			14'b01100100011101: M1r = 2'b00;
			14'b10100100011101: M1r = 2'b00;
			14'b11100100011101: M1r = 2'b00;
			14'b00110100011101: M1r = 2'b00;
			14'b01110100011101: M1r = 2'b00;
			14'b10110100011101: M1r = 2'b00;
			14'b11110100011101: M1r = 2'b00;
			14'b00001000011101: M1r = 2'b00;
			14'b01001000011101: M1r = 2'b00;
			14'b10001000011101: M1r = 2'b00;
			14'b11001000011101: M1r = 2'b00;
			14'b00011000011101: M1r = 2'b00;
			14'b01011000011101: M1r = 2'b00;
			14'b10011000011101: M1r = 2'b00;
			14'b11011000011101: M1r = 2'b00;
			14'b00101000011101: M1r = 2'b00;
			14'b01101000011101: M1r = 2'b00;
			14'b10101000011101: M1r = 2'b00;
			14'b11101000011101: M1r = 2'b00;
			14'b00111000011101: M1r = 2'b00;
			14'b01111000011101: M1r = 2'b00;
			14'b10111000011101: M1r = 2'b00;
			14'b11111000011101: M1r = 2'b00;
			14'b00001100011101: M1r = 2'b00;
			14'b01001100011101: M1r = 2'b01;
			14'b10001100011101: M1r = 2'b01;
			14'b11001100011101: M1r = 2'b01;
			14'b00011100011101: M1r = 2'b00;
			14'b01011100011101: M1r = 2'b00;
			14'b10011100011101: M1r = 2'b00;
			14'b11011100011101: M1r = 2'b00;
			14'b00101100011101: M1r = 2'b00;
			14'b01101100011101: M1r = 2'b00;
			14'b10101100011101: M1r = 2'b00;
			14'b11101100011101: M1r = 2'b00;
			14'b00111100011101: M1r = 2'b00;
			14'b01111100011101: M1r = 2'b00;
			14'b10111100011101: M1r = 2'b00;
			14'b11111100011101: M1r = 2'b00;
			14'b00000001011101: M1r = 2'b00;
			14'b01000001011101: M1r = 2'b00;
			14'b10000001011101: M1r = 2'b00;
			14'b11000001011101: M1r = 2'b00;
			14'b00010001011101: M1r = 2'b00;
			14'b01010001011101: M1r = 2'b00;
			14'b10010001011101: M1r = 2'b00;
			14'b11010001011101: M1r = 2'b00;
			14'b00100001011101: M1r = 2'b00;
			14'b01100001011101: M1r = 2'b00;
			14'b10100001011101: M1r = 2'b00;
			14'b11100001011101: M1r = 2'b00;
			14'b00110001011101: M1r = 2'b00;
			14'b01110001011101: M1r = 2'b00;
			14'b10110001011101: M1r = 2'b00;
			14'b11110001011101: M1r = 2'b00;
			14'b00000101011101: M1r = 2'b00;
			14'b01000101011101: M1r = 2'b00;
			14'b10000101011101: M1r = 2'b00;
			14'b11000101011101: M1r = 2'b00;
			14'b00010101011101: M1r = 2'b00;
			14'b01010101011101: M1r = 2'b00;
			14'b10010101011101: M1r = 2'b00;
			14'b11010101011101: M1r = 2'b00;
			14'b00100101011101: M1r = 2'b00;
			14'b01100101011101: M1r = 2'b00;
			14'b10100101011101: M1r = 2'b00;
			14'b11100101011101: M1r = 2'b00;
			14'b00110101011101: M1r = 2'b00;
			14'b01110101011101: M1r = 2'b00;
			14'b10110101011101: M1r = 2'b00;
			14'b11110101011101: M1r = 2'b00;
			14'b00001001011101: M1r = 2'b00;
			14'b01001001011101: M1r = 2'b00;
			14'b10001001011101: M1r = 2'b00;
			14'b11001001011101: M1r = 2'b00;
			14'b00011001011101: M1r = 2'b00;
			14'b01011001011101: M1r = 2'b00;
			14'b10011001011101: M1r = 2'b00;
			14'b11011001011101: M1r = 2'b00;
			14'b00101001011101: M1r = 2'b00;
			14'b01101001011101: M1r = 2'b00;
			14'b10101001011101: M1r = 2'b00;
			14'b11101001011101: M1r = 2'b00;
			14'b00111001011101: M1r = 2'b00;
			14'b01111001011101: M1r = 2'b00;
			14'b10111001011101: M1r = 2'b00;
			14'b11111001011101: M1r = 2'b00;
			14'b00001101011101: M1r = 2'b00;
			14'b01001101011101: M1r = 2'b00;
			14'b10001101011101: M1r = 2'b00;
			14'b11001101011101: M1r = 2'b01;
			14'b00011101011101: M1r = 2'b00;
			14'b01011101011101: M1r = 2'b00;
			14'b10011101011101: M1r = 2'b00;
			14'b11011101011101: M1r = 2'b00;
			14'b00101101011101: M1r = 2'b00;
			14'b01101101011101: M1r = 2'b00;
			14'b10101101011101: M1r = 2'b00;
			14'b11101101011101: M1r = 2'b00;
			14'b00111101011101: M1r = 2'b00;
			14'b01111101011101: M1r = 2'b00;
			14'b10111101011101: M1r = 2'b00;
			14'b11111101011101: M1r = 2'b00;
			14'b00000010011101: M1r = 2'b00;
			14'b01000010011101: M1r = 2'b00;
			14'b10000010011101: M1r = 2'b00;
			14'b11000010011101: M1r = 2'b00;
			14'b00010010011101: M1r = 2'b00;
			14'b01010010011101: M1r = 2'b00;
			14'b10010010011101: M1r = 2'b00;
			14'b11010010011101: M1r = 2'b00;
			14'b00100010011101: M1r = 2'b00;
			14'b01100010011101: M1r = 2'b00;
			14'b10100010011101: M1r = 2'b00;
			14'b11100010011101: M1r = 2'b00;
			14'b00110010011101: M1r = 2'b00;
			14'b01110010011101: M1r = 2'b00;
			14'b10110010011101: M1r = 2'b00;
			14'b11110010011101: M1r = 2'b00;
			14'b00000110011101: M1r = 2'b00;
			14'b01000110011101: M1r = 2'b00;
			14'b10000110011101: M1r = 2'b00;
			14'b11000110011101: M1r = 2'b00;
			14'b00010110011101: M1r = 2'b00;
			14'b01010110011101: M1r = 2'b00;
			14'b10010110011101: M1r = 2'b00;
			14'b11010110011101: M1r = 2'b00;
			14'b00100110011101: M1r = 2'b00;
			14'b01100110011101: M1r = 2'b00;
			14'b10100110011101: M1r = 2'b00;
			14'b11100110011101: M1r = 2'b00;
			14'b00110110011101: M1r = 2'b00;
			14'b01110110011101: M1r = 2'b00;
			14'b10110110011101: M1r = 2'b00;
			14'b11110110011101: M1r = 2'b00;
			14'b00001010011101: M1r = 2'b00;
			14'b01001010011101: M1r = 2'b00;
			14'b10001010011101: M1r = 2'b00;
			14'b11001010011101: M1r = 2'b00;
			14'b00011010011101: M1r = 2'b00;
			14'b01011010011101: M1r = 2'b00;
			14'b10011010011101: M1r = 2'b00;
			14'b11011010011101: M1r = 2'b00;
			14'b00101010011101: M1r = 2'b00;
			14'b01101010011101: M1r = 2'b00;
			14'b10101010011101: M1r = 2'b00;
			14'b11101010011101: M1r = 2'b00;
			14'b00111010011101: M1r = 2'b00;
			14'b01111010011101: M1r = 2'b00;
			14'b10111010011101: M1r = 2'b00;
			14'b11111010011101: M1r = 2'b00;
			14'b00001110011101: M1r = 2'b00;
			14'b01001110011101: M1r = 2'b00;
			14'b10001110011101: M1r = 2'b00;
			14'b11001110011101: M1r = 2'b00;
			14'b00011110011101: M1r = 2'b00;
			14'b01011110011101: M1r = 2'b00;
			14'b10011110011101: M1r = 2'b00;
			14'b11011110011101: M1r = 2'b00;
			14'b00101110011101: M1r = 2'b00;
			14'b01101110011101: M1r = 2'b00;
			14'b10101110011101: M1r = 2'b00;
			14'b11101110011101: M1r = 2'b00;
			14'b00111110011101: M1r = 2'b00;
			14'b01111110011101: M1r = 2'b00;
			14'b10111110011101: M1r = 2'b00;
			14'b11111110011101: M1r = 2'b00;
			14'b00000011011101: M1r = 2'b00;
			14'b01000011011101: M1r = 2'b00;
			14'b10000011011101: M1r = 2'b00;
			14'b11000011011101: M1r = 2'b00;
			14'b00010011011101: M1r = 2'b00;
			14'b01010011011101: M1r = 2'b00;
			14'b10010011011101: M1r = 2'b00;
			14'b11010011011101: M1r = 2'b00;
			14'b00100011011101: M1r = 2'b00;
			14'b01100011011101: M1r = 2'b00;
			14'b10100011011101: M1r = 2'b00;
			14'b11100011011101: M1r = 2'b00;
			14'b00110011011101: M1r = 2'b00;
			14'b01110011011101: M1r = 2'b00;
			14'b10110011011101: M1r = 2'b00;
			14'b11110011011101: M1r = 2'b00;
			14'b00000111011101: M1r = 2'b00;
			14'b01000111011101: M1r = 2'b00;
			14'b10000111011101: M1r = 2'b00;
			14'b11000111011101: M1r = 2'b00;
			14'b00010111011101: M1r = 2'b00;
			14'b01010111011101: M1r = 2'b00;
			14'b10010111011101: M1r = 2'b00;
			14'b11010111011101: M1r = 2'b00;
			14'b00100111011101: M1r = 2'b00;
			14'b01100111011101: M1r = 2'b00;
			14'b10100111011101: M1r = 2'b00;
			14'b11100111011101: M1r = 2'b00;
			14'b00110111011101: M1r = 2'b00;
			14'b01110111011101: M1r = 2'b00;
			14'b10110111011101: M1r = 2'b00;
			14'b11110111011101: M1r = 2'b00;
			14'b00001011011101: M1r = 2'b00;
			14'b01001011011101: M1r = 2'b00;
			14'b10001011011101: M1r = 2'b00;
			14'b11001011011101: M1r = 2'b00;
			14'b00011011011101: M1r = 2'b00;
			14'b01011011011101: M1r = 2'b00;
			14'b10011011011101: M1r = 2'b00;
			14'b11011011011101: M1r = 2'b00;
			14'b00101011011101: M1r = 2'b00;
			14'b01101011011101: M1r = 2'b00;
			14'b10101011011101: M1r = 2'b00;
			14'b11101011011101: M1r = 2'b00;
			14'b00111011011101: M1r = 2'b00;
			14'b01111011011101: M1r = 2'b00;
			14'b10111011011101: M1r = 2'b00;
			14'b11111011011101: M1r = 2'b00;
			14'b00001111011101: M1r = 2'b00;
			14'b01001111011101: M1r = 2'b00;
			14'b10001111011101: M1r = 2'b00;
			14'b11001111011101: M1r = 2'b00;
			14'b00011111011101: M1r = 2'b00;
			14'b01011111011101: M1r = 2'b00;
			14'b10011111011101: M1r = 2'b00;
			14'b11011111011101: M1r = 2'b00;
			14'b00101111011101: M1r = 2'b00;
			14'b01101111011101: M1r = 2'b00;
			14'b10101111011101: M1r = 2'b00;
			14'b11101111011101: M1r = 2'b00;
			14'b00111111011101: M1r = 2'b00;
			14'b01111111011101: M1r = 2'b00;
			14'b10111111011101: M1r = 2'b00;
			14'b11111111011101: M1r = 2'b00;
			14'b00000000101101: M1r = 2'b00;
			14'b01000000101101: M1r = 2'b00;
			14'b10000000101101: M1r = 2'b00;
			14'b11000000101101: M1r = 2'b00;
			14'b00010000101101: M1r = 2'b00;
			14'b01010000101101: M1r = 2'b00;
			14'b10010000101101: M1r = 2'b00;
			14'b11010000101101: M1r = 2'b00;
			14'b00100000101101: M1r = 2'b00;
			14'b01100000101101: M1r = 2'b00;
			14'b10100000101101: M1r = 2'b00;
			14'b11100000101101: M1r = 2'b00;
			14'b00110000101101: M1r = 2'b00;
			14'b01110000101101: M1r = 2'b00;
			14'b10110000101101: M1r = 2'b00;
			14'b11110000101101: M1r = 2'b00;
			14'b00000100101101: M1r = 2'b00;
			14'b01000100101101: M1r = 2'b00;
			14'b10000100101101: M1r = 2'b00;
			14'b11000100101101: M1r = 2'b00;
			14'b00010100101101: M1r = 2'b00;
			14'b01010100101101: M1r = 2'b00;
			14'b10010100101101: M1r = 2'b00;
			14'b11010100101101: M1r = 2'b00;
			14'b00100100101101: M1r = 2'b00;
			14'b01100100101101: M1r = 2'b00;
			14'b10100100101101: M1r = 2'b00;
			14'b11100100101101: M1r = 2'b00;
			14'b00110100101101: M1r = 2'b00;
			14'b01110100101101: M1r = 2'b00;
			14'b10110100101101: M1r = 2'b00;
			14'b11110100101101: M1r = 2'b00;
			14'b00001000101101: M1r = 2'b00;
			14'b01001000101101: M1r = 2'b00;
			14'b10001000101101: M1r = 2'b00;
			14'b11001000101101: M1r = 2'b01;
			14'b00011000101101: M1r = 2'b00;
			14'b01011000101101: M1r = 2'b00;
			14'b10011000101101: M1r = 2'b00;
			14'b11011000101101: M1r = 2'b00;
			14'b00101000101101: M1r = 2'b00;
			14'b01101000101101: M1r = 2'b00;
			14'b10101000101101: M1r = 2'b00;
			14'b11101000101101: M1r = 2'b00;
			14'b00111000101101: M1r = 2'b00;
			14'b01111000101101: M1r = 2'b00;
			14'b10111000101101: M1r = 2'b00;
			14'b11111000101101: M1r = 2'b00;
			14'b00001100101101: M1r = 2'b01;
			14'b01001100101101: M1r = 2'b01;
			14'b10001100101101: M1r = 2'b01;
			14'b11001100101101: M1r = 2'b01;
			14'b00011100101101: M1r = 2'b00;
			14'b01011100101101: M1r = 2'b01;
			14'b10011100101101: M1r = 2'b01;
			14'b11011100101101: M1r = 2'b01;
			14'b00101100101101: M1r = 2'b00;
			14'b01101100101101: M1r = 2'b00;
			14'b10101100101101: M1r = 2'b00;
			14'b11101100101101: M1r = 2'b00;
			14'b00111100101101: M1r = 2'b00;
			14'b01111100101101: M1r = 2'b00;
			14'b10111100101101: M1r = 2'b00;
			14'b11111100101101: M1r = 2'b00;
			14'b00000001101101: M1r = 2'b00;
			14'b01000001101101: M1r = 2'b00;
			14'b10000001101101: M1r = 2'b00;
			14'b11000001101101: M1r = 2'b00;
			14'b00010001101101: M1r = 2'b00;
			14'b01010001101101: M1r = 2'b00;
			14'b10010001101101: M1r = 2'b00;
			14'b11010001101101: M1r = 2'b00;
			14'b00100001101101: M1r = 2'b00;
			14'b01100001101101: M1r = 2'b00;
			14'b10100001101101: M1r = 2'b00;
			14'b11100001101101: M1r = 2'b00;
			14'b00110001101101: M1r = 2'b00;
			14'b01110001101101: M1r = 2'b00;
			14'b10110001101101: M1r = 2'b00;
			14'b11110001101101: M1r = 2'b00;
			14'b00000101101101: M1r = 2'b00;
			14'b01000101101101: M1r = 2'b00;
			14'b10000101101101: M1r = 2'b00;
			14'b11000101101101: M1r = 2'b00;
			14'b00010101101101: M1r = 2'b00;
			14'b01010101101101: M1r = 2'b00;
			14'b10010101101101: M1r = 2'b00;
			14'b11010101101101: M1r = 2'b00;
			14'b00100101101101: M1r = 2'b00;
			14'b01100101101101: M1r = 2'b00;
			14'b10100101101101: M1r = 2'b00;
			14'b11100101101101: M1r = 2'b00;
			14'b00110101101101: M1r = 2'b00;
			14'b01110101101101: M1r = 2'b00;
			14'b10110101101101: M1r = 2'b00;
			14'b11110101101101: M1r = 2'b00;
			14'b00001001101101: M1r = 2'b00;
			14'b01001001101101: M1r = 2'b00;
			14'b10001001101101: M1r = 2'b00;
			14'b11001001101101: M1r = 2'b00;
			14'b00011001101101: M1r = 2'b00;
			14'b01011001101101: M1r = 2'b00;
			14'b10011001101101: M1r = 2'b00;
			14'b11011001101101: M1r = 2'b00;
			14'b00101001101101: M1r = 2'b00;
			14'b01101001101101: M1r = 2'b00;
			14'b10101001101101: M1r = 2'b00;
			14'b11101001101101: M1r = 2'b00;
			14'b00111001101101: M1r = 2'b00;
			14'b01111001101101: M1r = 2'b00;
			14'b10111001101101: M1r = 2'b00;
			14'b11111001101101: M1r = 2'b00;
			14'b00001101101101: M1r = 2'b01;
			14'b01001101101101: M1r = 2'b01;
			14'b10001101101101: M1r = 2'b01;
			14'b11001101101101: M1r = 2'b01;
			14'b00011101101101: M1r = 2'b00;
			14'b01011101101101: M1r = 2'b00;
			14'b10011101101101: M1r = 2'b00;
			14'b11011101101101: M1r = 2'b01;
			14'b00101101101101: M1r = 2'b00;
			14'b01101101101101: M1r = 2'b00;
			14'b10101101101101: M1r = 2'b00;
			14'b11101101101101: M1r = 2'b00;
			14'b00111101101101: M1r = 2'b00;
			14'b01111101101101: M1r = 2'b00;
			14'b10111101101101: M1r = 2'b00;
			14'b11111101101101: M1r = 2'b00;
			14'b00000010101101: M1r = 2'b00;
			14'b01000010101101: M1r = 2'b00;
			14'b10000010101101: M1r = 2'b00;
			14'b11000010101101: M1r = 2'b00;
			14'b00010010101101: M1r = 2'b00;
			14'b01010010101101: M1r = 2'b00;
			14'b10010010101101: M1r = 2'b00;
			14'b11010010101101: M1r = 2'b00;
			14'b00100010101101: M1r = 2'b00;
			14'b01100010101101: M1r = 2'b00;
			14'b10100010101101: M1r = 2'b00;
			14'b11100010101101: M1r = 2'b00;
			14'b00110010101101: M1r = 2'b00;
			14'b01110010101101: M1r = 2'b00;
			14'b10110010101101: M1r = 2'b00;
			14'b11110010101101: M1r = 2'b00;
			14'b00000110101101: M1r = 2'b00;
			14'b01000110101101: M1r = 2'b00;
			14'b10000110101101: M1r = 2'b00;
			14'b11000110101101: M1r = 2'b00;
			14'b00010110101101: M1r = 2'b00;
			14'b01010110101101: M1r = 2'b00;
			14'b10010110101101: M1r = 2'b00;
			14'b11010110101101: M1r = 2'b00;
			14'b00100110101101: M1r = 2'b00;
			14'b01100110101101: M1r = 2'b00;
			14'b10100110101101: M1r = 2'b00;
			14'b11100110101101: M1r = 2'b00;
			14'b00110110101101: M1r = 2'b00;
			14'b01110110101101: M1r = 2'b00;
			14'b10110110101101: M1r = 2'b00;
			14'b11110110101101: M1r = 2'b00;
			14'b00001010101101: M1r = 2'b00;
			14'b01001010101101: M1r = 2'b00;
			14'b10001010101101: M1r = 2'b00;
			14'b11001010101101: M1r = 2'b00;
			14'b00011010101101: M1r = 2'b00;
			14'b01011010101101: M1r = 2'b00;
			14'b10011010101101: M1r = 2'b00;
			14'b11011010101101: M1r = 2'b00;
			14'b00101010101101: M1r = 2'b00;
			14'b01101010101101: M1r = 2'b00;
			14'b10101010101101: M1r = 2'b00;
			14'b11101010101101: M1r = 2'b00;
			14'b00111010101101: M1r = 2'b00;
			14'b01111010101101: M1r = 2'b00;
			14'b10111010101101: M1r = 2'b00;
			14'b11111010101101: M1r = 2'b00;
			14'b00001110101101: M1r = 2'b00;
			14'b01001110101101: M1r = 2'b00;
			14'b10001110101101: M1r = 2'b01;
			14'b11001110101101: M1r = 2'b01;
			14'b00011110101101: M1r = 2'b00;
			14'b01011110101101: M1r = 2'b00;
			14'b10011110101101: M1r = 2'b00;
			14'b11011110101101: M1r = 2'b00;
			14'b00101110101101: M1r = 2'b00;
			14'b01101110101101: M1r = 2'b00;
			14'b10101110101101: M1r = 2'b00;
			14'b11101110101101: M1r = 2'b00;
			14'b00111110101101: M1r = 2'b00;
			14'b01111110101101: M1r = 2'b00;
			14'b10111110101101: M1r = 2'b00;
			14'b11111110101101: M1r = 2'b00;
			14'b00000011101101: M1r = 2'b00;
			14'b01000011101101: M1r = 2'b00;
			14'b10000011101101: M1r = 2'b00;
			14'b11000011101101: M1r = 2'b00;
			14'b00010011101101: M1r = 2'b00;
			14'b01010011101101: M1r = 2'b00;
			14'b10010011101101: M1r = 2'b00;
			14'b11010011101101: M1r = 2'b00;
			14'b00100011101101: M1r = 2'b00;
			14'b01100011101101: M1r = 2'b00;
			14'b10100011101101: M1r = 2'b00;
			14'b11100011101101: M1r = 2'b00;
			14'b00110011101101: M1r = 2'b00;
			14'b01110011101101: M1r = 2'b00;
			14'b10110011101101: M1r = 2'b00;
			14'b11110011101101: M1r = 2'b00;
			14'b00000111101101: M1r = 2'b00;
			14'b01000111101101: M1r = 2'b00;
			14'b10000111101101: M1r = 2'b00;
			14'b11000111101101: M1r = 2'b00;
			14'b00010111101101: M1r = 2'b00;
			14'b01010111101101: M1r = 2'b00;
			14'b10010111101101: M1r = 2'b00;
			14'b11010111101101: M1r = 2'b00;
			14'b00100111101101: M1r = 2'b00;
			14'b01100111101101: M1r = 2'b00;
			14'b10100111101101: M1r = 2'b00;
			14'b11100111101101: M1r = 2'b00;
			14'b00110111101101: M1r = 2'b00;
			14'b01110111101101: M1r = 2'b00;
			14'b10110111101101: M1r = 2'b00;
			14'b11110111101101: M1r = 2'b00;
			14'b00001011101101: M1r = 2'b00;
			14'b01001011101101: M1r = 2'b00;
			14'b10001011101101: M1r = 2'b00;
			14'b11001011101101: M1r = 2'b00;
			14'b00011011101101: M1r = 2'b00;
			14'b01011011101101: M1r = 2'b00;
			14'b10011011101101: M1r = 2'b00;
			14'b11011011101101: M1r = 2'b00;
			14'b00101011101101: M1r = 2'b00;
			14'b01101011101101: M1r = 2'b00;
			14'b10101011101101: M1r = 2'b00;
			14'b11101011101101: M1r = 2'b00;
			14'b00111011101101: M1r = 2'b00;
			14'b01111011101101: M1r = 2'b00;
			14'b10111011101101: M1r = 2'b00;
			14'b11111011101101: M1r = 2'b00;
			14'b00001111101101: M1r = 2'b00;
			14'b01001111101101: M1r = 2'b00;
			14'b10001111101101: M1r = 2'b00;
			14'b11001111101101: M1r = 2'b01;
			14'b00011111101101: M1r = 2'b00;
			14'b01011111101101: M1r = 2'b00;
			14'b10011111101101: M1r = 2'b00;
			14'b11011111101101: M1r = 2'b00;
			14'b00101111101101: M1r = 2'b00;
			14'b01101111101101: M1r = 2'b00;
			14'b10101111101101: M1r = 2'b00;
			14'b11101111101101: M1r = 2'b00;
			14'b00111111101101: M1r = 2'b00;
			14'b01111111101101: M1r = 2'b00;
			14'b10111111101101: M1r = 2'b00;
			14'b11111111101101: M1r = 2'b00;
			14'b00000000111101: M1r = 2'b00;
			14'b01000000111101: M1r = 2'b00;
			14'b10000000111101: M1r = 2'b00;
			14'b11000000111101: M1r = 2'b00;
			14'b00010000111101: M1r = 2'b00;
			14'b01010000111101: M1r = 2'b00;
			14'b10010000111101: M1r = 2'b00;
			14'b11010000111101: M1r = 2'b00;
			14'b00100000111101: M1r = 2'b00;
			14'b01100000111101: M1r = 2'b00;
			14'b10100000111101: M1r = 2'b00;
			14'b11100000111101: M1r = 2'b00;
			14'b00110000111101: M1r = 2'b00;
			14'b01110000111101: M1r = 2'b00;
			14'b10110000111101: M1r = 2'b00;
			14'b11110000111101: M1r = 2'b00;
			14'b00000100111101: M1r = 2'b00;
			14'b01000100111101: M1r = 2'b00;
			14'b10000100111101: M1r = 2'b00;
			14'b11000100111101: M1r = 2'b00;
			14'b00010100111101: M1r = 2'b00;
			14'b01010100111101: M1r = 2'b00;
			14'b10010100111101: M1r = 2'b00;
			14'b11010100111101: M1r = 2'b00;
			14'b00100100111101: M1r = 2'b00;
			14'b01100100111101: M1r = 2'b00;
			14'b10100100111101: M1r = 2'b00;
			14'b11100100111101: M1r = 2'b00;
			14'b00110100111101: M1r = 2'b00;
			14'b01110100111101: M1r = 2'b00;
			14'b10110100111101: M1r = 2'b00;
			14'b11110100111101: M1r = 2'b00;
			14'b00001000111101: M1r = 2'b01;
			14'b01001000111101: M1r = 2'b01;
			14'b10001000111101: M1r = 2'b01;
			14'b11001000111101: M1r = 2'b01;
			14'b00011000111101: M1r = 2'b00;
			14'b01011000111101: M1r = 2'b00;
			14'b10011000111101: M1r = 2'b00;
			14'b11011000111101: M1r = 2'b01;
			14'b00101000111101: M1r = 2'b00;
			14'b01101000111101: M1r = 2'b00;
			14'b10101000111101: M1r = 2'b00;
			14'b11101000111101: M1r = 2'b00;
			14'b00111000111101: M1r = 2'b00;
			14'b01111000111101: M1r = 2'b00;
			14'b10111000111101: M1r = 2'b00;
			14'b11111000111101: M1r = 2'b00;
			14'b00001100111101: M1r = 2'b01;
			14'b01001100111101: M1r = 2'b01;
			14'b10001100111101: M1r = 2'b10;
			14'b11001100111101: M1r = 2'b10;
			14'b00011100111101: M1r = 2'b01;
			14'b01011100111101: M1r = 2'b01;
			14'b10011100111101: M1r = 2'b01;
			14'b11011100111101: M1r = 2'b01;
			14'b00101100111101: M1r = 2'b00;
			14'b01101100111101: M1r = 2'b01;
			14'b10101100111101: M1r = 2'b01;
			14'b11101100111101: M1r = 2'b01;
			14'b00111100111101: M1r = 2'b00;
			14'b01111100111101: M1r = 2'b00;
			14'b10111100111101: M1r = 2'b00;
			14'b11111100111101: M1r = 2'b00;
			14'b00000001111101: M1r = 2'b00;
			14'b01000001111101: M1r = 2'b00;
			14'b10000001111101: M1r = 2'b00;
			14'b11000001111101: M1r = 2'b00;
			14'b00010001111101: M1r = 2'b00;
			14'b01010001111101: M1r = 2'b00;
			14'b10010001111101: M1r = 2'b00;
			14'b11010001111101: M1r = 2'b00;
			14'b00100001111101: M1r = 2'b00;
			14'b01100001111101: M1r = 2'b00;
			14'b10100001111101: M1r = 2'b00;
			14'b11100001111101: M1r = 2'b00;
			14'b00110001111101: M1r = 2'b00;
			14'b01110001111101: M1r = 2'b00;
			14'b10110001111101: M1r = 2'b00;
			14'b11110001111101: M1r = 2'b00;
			14'b00000101111101: M1r = 2'b00;
			14'b01000101111101: M1r = 2'b00;
			14'b10000101111101: M1r = 2'b00;
			14'b11000101111101: M1r = 2'b00;
			14'b00010101111101: M1r = 2'b00;
			14'b01010101111101: M1r = 2'b00;
			14'b10010101111101: M1r = 2'b00;
			14'b11010101111101: M1r = 2'b00;
			14'b00100101111101: M1r = 2'b00;
			14'b01100101111101: M1r = 2'b00;
			14'b10100101111101: M1r = 2'b00;
			14'b11100101111101: M1r = 2'b00;
			14'b00110101111101: M1r = 2'b00;
			14'b01110101111101: M1r = 2'b00;
			14'b10110101111101: M1r = 2'b00;
			14'b11110101111101: M1r = 2'b00;
			14'b00001001111101: M1r = 2'b00;
			14'b01001001111101: M1r = 2'b00;
			14'b10001001111101: M1r = 2'b01;
			14'b11001001111101: M1r = 2'b01;
			14'b00011001111101: M1r = 2'b00;
			14'b01011001111101: M1r = 2'b00;
			14'b10011001111101: M1r = 2'b00;
			14'b11011001111101: M1r = 2'b00;
			14'b00101001111101: M1r = 2'b00;
			14'b01101001111101: M1r = 2'b00;
			14'b10101001111101: M1r = 2'b00;
			14'b11101001111101: M1r = 2'b00;
			14'b00111001111101: M1r = 2'b00;
			14'b01111001111101: M1r = 2'b00;
			14'b10111001111101: M1r = 2'b00;
			14'b11111001111101: M1r = 2'b00;
			14'b00001101111101: M1r = 2'b01;
			14'b01001101111101: M1r = 2'b01;
			14'b10001101111101: M1r = 2'b01;
			14'b11001101111101: M1r = 2'b10;
			14'b00011101111101: M1r = 2'b01;
			14'b01011101111101: M1r = 2'b01;
			14'b10011101111101: M1r = 2'b01;
			14'b11011101111101: M1r = 2'b01;
			14'b00101101111101: M1r = 2'b00;
			14'b01101101111101: M1r = 2'b00;
			14'b10101101111101: M1r = 2'b00;
			14'b11101101111101: M1r = 2'b01;
			14'b00111101111101: M1r = 2'b00;
			14'b01111101111101: M1r = 2'b00;
			14'b10111101111101: M1r = 2'b00;
			14'b11111101111101: M1r = 2'b00;
			14'b00000010111101: M1r = 2'b00;
			14'b01000010111101: M1r = 2'b00;
			14'b10000010111101: M1r = 2'b00;
			14'b11000010111101: M1r = 2'b00;
			14'b00010010111101: M1r = 2'b00;
			14'b01010010111101: M1r = 2'b00;
			14'b10010010111101: M1r = 2'b00;
			14'b11010010111101: M1r = 2'b00;
			14'b00100010111101: M1r = 2'b00;
			14'b01100010111101: M1r = 2'b00;
			14'b10100010111101: M1r = 2'b00;
			14'b11100010111101: M1r = 2'b00;
			14'b00110010111101: M1r = 2'b00;
			14'b01110010111101: M1r = 2'b00;
			14'b10110010111101: M1r = 2'b00;
			14'b11110010111101: M1r = 2'b00;
			14'b00000110111101: M1r = 2'b00;
			14'b01000110111101: M1r = 2'b00;
			14'b10000110111101: M1r = 2'b00;
			14'b11000110111101: M1r = 2'b00;
			14'b00010110111101: M1r = 2'b00;
			14'b01010110111101: M1r = 2'b00;
			14'b10010110111101: M1r = 2'b00;
			14'b11010110111101: M1r = 2'b00;
			14'b00100110111101: M1r = 2'b00;
			14'b01100110111101: M1r = 2'b00;
			14'b10100110111101: M1r = 2'b00;
			14'b11100110111101: M1r = 2'b00;
			14'b00110110111101: M1r = 2'b00;
			14'b01110110111101: M1r = 2'b00;
			14'b10110110111101: M1r = 2'b00;
			14'b11110110111101: M1r = 2'b00;
			14'b00001010111101: M1r = 2'b00;
			14'b01001010111101: M1r = 2'b00;
			14'b10001010111101: M1r = 2'b00;
			14'b11001010111101: M1r = 2'b00;
			14'b00011010111101: M1r = 2'b00;
			14'b01011010111101: M1r = 2'b00;
			14'b10011010111101: M1r = 2'b00;
			14'b11011010111101: M1r = 2'b00;
			14'b00101010111101: M1r = 2'b00;
			14'b01101010111101: M1r = 2'b00;
			14'b10101010111101: M1r = 2'b00;
			14'b11101010111101: M1r = 2'b00;
			14'b00111010111101: M1r = 2'b00;
			14'b01111010111101: M1r = 2'b00;
			14'b10111010111101: M1r = 2'b00;
			14'b11111010111101: M1r = 2'b00;
			14'b00001110111101: M1r = 2'b01;
			14'b01001110111101: M1r = 2'b01;
			14'b10001110111101: M1r = 2'b01;
			14'b11001110111101: M1r = 2'b01;
			14'b00011110111101: M1r = 2'b00;
			14'b01011110111101: M1r = 2'b00;
			14'b10011110111101: M1r = 2'b01;
			14'b11011110111101: M1r = 2'b01;
			14'b00101110111101: M1r = 2'b00;
			14'b01101110111101: M1r = 2'b00;
			14'b10101110111101: M1r = 2'b00;
			14'b11101110111101: M1r = 2'b00;
			14'b00111110111101: M1r = 2'b00;
			14'b01111110111101: M1r = 2'b00;
			14'b10111110111101: M1r = 2'b00;
			14'b11111110111101: M1r = 2'b00;
			14'b00000011111101: M1r = 2'b00;
			14'b01000011111101: M1r = 2'b00;
			14'b10000011111101: M1r = 2'b00;
			14'b11000011111101: M1r = 2'b00;
			14'b00010011111101: M1r = 2'b00;
			14'b01010011111101: M1r = 2'b00;
			14'b10010011111101: M1r = 2'b00;
			14'b11010011111101: M1r = 2'b00;
			14'b00100011111101: M1r = 2'b00;
			14'b01100011111101: M1r = 2'b00;
			14'b10100011111101: M1r = 2'b00;
			14'b11100011111101: M1r = 2'b00;
			14'b00110011111101: M1r = 2'b00;
			14'b01110011111101: M1r = 2'b00;
			14'b10110011111101: M1r = 2'b00;
			14'b11110011111101: M1r = 2'b00;
			14'b00000111111101: M1r = 2'b00;
			14'b01000111111101: M1r = 2'b00;
			14'b10000111111101: M1r = 2'b00;
			14'b11000111111101: M1r = 2'b00;
			14'b00010111111101: M1r = 2'b00;
			14'b01010111111101: M1r = 2'b00;
			14'b10010111111101: M1r = 2'b00;
			14'b11010111111101: M1r = 2'b00;
			14'b00100111111101: M1r = 2'b00;
			14'b01100111111101: M1r = 2'b00;
			14'b10100111111101: M1r = 2'b00;
			14'b11100111111101: M1r = 2'b00;
			14'b00110111111101: M1r = 2'b00;
			14'b01110111111101: M1r = 2'b00;
			14'b10110111111101: M1r = 2'b00;
			14'b11110111111101: M1r = 2'b00;
			14'b00001011111101: M1r = 2'b00;
			14'b01001011111101: M1r = 2'b00;
			14'b10001011111101: M1r = 2'b00;
			14'b11001011111101: M1r = 2'b00;
			14'b00011011111101: M1r = 2'b00;
			14'b01011011111101: M1r = 2'b00;
			14'b10011011111101: M1r = 2'b00;
			14'b11011011111101: M1r = 2'b00;
			14'b00101011111101: M1r = 2'b00;
			14'b01101011111101: M1r = 2'b00;
			14'b10101011111101: M1r = 2'b00;
			14'b11101011111101: M1r = 2'b00;
			14'b00111011111101: M1r = 2'b00;
			14'b01111011111101: M1r = 2'b00;
			14'b10111011111101: M1r = 2'b00;
			14'b11111011111101: M1r = 2'b00;
			14'b00001111111101: M1r = 2'b00;
			14'b01001111111101: M1r = 2'b01;
			14'b10001111111101: M1r = 2'b01;
			14'b11001111111101: M1r = 2'b01;
			14'b00011111111101: M1r = 2'b00;
			14'b01011111111101: M1r = 2'b00;
			14'b10011111111101: M1r = 2'b00;
			14'b11011111111101: M1r = 2'b00;
			14'b00101111111101: M1r = 2'b00;
			14'b01101111111101: M1r = 2'b00;
			14'b10101111111101: M1r = 2'b00;
			14'b11101111111101: M1r = 2'b00;
			14'b00111111111101: M1r = 2'b00;
			14'b01111111111101: M1r = 2'b00;
			14'b10111111111101: M1r = 2'b00;
			14'b11111111111101: M1r = 2'b00;
			14'b00000000000010: M1r = 2'b01;
			14'b01000000000010: M1r = 2'b01;
			14'b10000000000010: M1r = 2'b01;
			14'b11000000000010: M1r = 2'b10;
			14'b00010000000010: M1r = 2'b01;
			14'b01010000000010: M1r = 2'b01;
			14'b10010000000010: M1r = 2'b01;
			14'b11010000000010: M1r = 2'b01;
			14'b00100000000010: M1r = 2'b00;
			14'b01100000000010: M1r = 2'b00;
			14'b10100000000010: M1r = 2'b00;
			14'b11100000000010: M1r = 2'b01;
			14'b00110000000010: M1r = 2'b00;
			14'b01110000000010: M1r = 2'b00;
			14'b10110000000010: M1r = 2'b00;
			14'b11110000000010: M1r = 2'b00;
			14'b00000100000010: M1r = 2'b10;
			14'b01000100000010: M1r = 2'b10;
			14'b10000100000010: M1r = 2'b10;
			14'b11000100000010: M1r = 2'b10;
			14'b00010100000010: M1r = 2'b01;
			14'b01010100000010: M1r = 2'b10;
			14'b10010100000010: M1r = 2'b10;
			14'b11010100000010: M1r = 2'b10;
			14'b00100100000010: M1r = 2'b01;
			14'b01100100000010: M1r = 2'b01;
			14'b10100100000010: M1r = 2'b01;
			14'b11100100000010: M1r = 2'b01;
			14'b00110100000010: M1r = 2'b00;
			14'b01110100000010: M1r = 2'b01;
			14'b10110100000010: M1r = 2'b01;
			14'b11110100000010: M1r = 2'b01;
			14'b00001000000010: M1r = 2'b11;
			14'b01001000000010: M1r = 2'b11;
			14'b10001000000010: M1r = 2'b11;
			14'b11001000000010: M1r = 2'b11;
			14'b00011000000010: M1r = 2'b10;
			14'b01011000000010: M1r = 2'b10;
			14'b10011000000010: M1r = 2'b10;
			14'b11011000000010: M1r = 2'b11;
			14'b00101000000010: M1r = 2'b10;
			14'b01101000000010: M1r = 2'b10;
			14'b10101000000010: M1r = 2'b10;
			14'b11101000000010: M1r = 2'b10;
			14'b00111000000010: M1r = 2'b01;
			14'b01111000000010: M1r = 2'b01;
			14'b10111000000010: M1r = 2'b01;
			14'b11111000000010: M1r = 2'b10;
			14'b00001100000010: M1r = 2'b11;
			14'b01001100000010: M1r = 2'b11;
			14'b10001100000010: M1r = 2'b11;
			14'b11001100000010: M1r = 2'b11;
			14'b00011100000010: M1r = 2'b11;
			14'b01011100000010: M1r = 2'b11;
			14'b10011100000010: M1r = 2'b11;
			14'b11011100000010: M1r = 2'b11;
			14'b00101100000010: M1r = 2'b10;
			14'b01101100000010: M1r = 2'b11;
			14'b10101100000010: M1r = 2'b11;
			14'b11101100000010: M1r = 2'b11;
			14'b00111100000010: M1r = 2'b10;
			14'b01111100000010: M1r = 2'b10;
			14'b10111100000010: M1r = 2'b10;
			14'b11111100000010: M1r = 2'b10;
			14'b00000001000010: M1r = 2'b01;
			14'b01000001000010: M1r = 2'b01;
			14'b10000001000010: M1r = 2'b01;
			14'b11000001000010: M1r = 2'b01;
			14'b00010001000010: M1r = 2'b00;
			14'b01010001000010: M1r = 2'b00;
			14'b10010001000010: M1r = 2'b01;
			14'b11010001000010: M1r = 2'b01;
			14'b00100001000010: M1r = 2'b00;
			14'b01100001000010: M1r = 2'b00;
			14'b10100001000010: M1r = 2'b00;
			14'b11100001000010: M1r = 2'b00;
			14'b00110001000010: M1r = 2'b00;
			14'b01110001000010: M1r = 2'b00;
			14'b10110001000010: M1r = 2'b00;
			14'b11110001000010: M1r = 2'b00;
			14'b00000101000010: M1r = 2'b10;
			14'b01000101000010: M1r = 2'b10;
			14'b10000101000010: M1r = 2'b10;
			14'b11000101000010: M1r = 2'b10;
			14'b00010101000010: M1r = 2'b01;
			14'b01010101000010: M1r = 2'b01;
			14'b10010101000010: M1r = 2'b01;
			14'b11010101000010: M1r = 2'b10;
			14'b00100101000010: M1r = 2'b01;
			14'b01100101000010: M1r = 2'b01;
			14'b10100101000010: M1r = 2'b01;
			14'b11100101000010: M1r = 2'b01;
			14'b00110101000010: M1r = 2'b00;
			14'b01110101000010: M1r = 2'b00;
			14'b10110101000010: M1r = 2'b00;
			14'b11110101000010: M1r = 2'b01;
			14'b00001001000010: M1r = 2'b10;
			14'b01001001000010: M1r = 2'b10;
			14'b10001001000010: M1r = 2'b11;
			14'b11001001000010: M1r = 2'b11;
			14'b00011001000010: M1r = 2'b10;
			14'b01011001000010: M1r = 2'b10;
			14'b10011001000010: M1r = 2'b10;
			14'b11011001000010: M1r = 2'b10;
			14'b00101001000010: M1r = 2'b01;
			14'b01101001000010: M1r = 2'b10;
			14'b10101001000010: M1r = 2'b10;
			14'b11101001000010: M1r = 2'b10;
			14'b00111001000010: M1r = 2'b01;
			14'b01111001000010: M1r = 2'b01;
			14'b10111001000010: M1r = 2'b01;
			14'b11111001000010: M1r = 2'b01;
			14'b00001101000010: M1r = 2'b11;
			14'b01001101000010: M1r = 2'b11;
			14'b10001101000010: M1r = 2'b11;
			14'b11001101000010: M1r = 2'b11;
			14'b00011101000010: M1r = 2'b11;
			14'b01011101000010: M1r = 2'b11;
			14'b10011101000010: M1r = 2'b11;
			14'b11011101000010: M1r = 2'b11;
			14'b00101101000010: M1r = 2'b10;
			14'b01101101000010: M1r = 2'b10;
			14'b10101101000010: M1r = 2'b10;
			14'b11101101000010: M1r = 2'b11;
			14'b00111101000010: M1r = 2'b10;
			14'b01111101000010: M1r = 2'b10;
			14'b10111101000010: M1r = 2'b10;
			14'b11111101000010: M1r = 2'b10;
			14'b00000010000010: M1r = 2'b01;
			14'b01000010000010: M1r = 2'b01;
			14'b10000010000010: M1r = 2'b01;
			14'b11000010000010: M1r = 2'b01;
			14'b00010010000010: M1r = 2'b00;
			14'b01010010000010: M1r = 2'b00;
			14'b10010010000010: M1r = 2'b00;
			14'b11010010000010: M1r = 2'b01;
			14'b00100010000010: M1r = 2'b00;
			14'b01100010000010: M1r = 2'b00;
			14'b10100010000010: M1r = 2'b00;
			14'b11100010000010: M1r = 2'b00;
			14'b00110010000010: M1r = 2'b00;
			14'b01110010000010: M1r = 2'b00;
			14'b10110010000010: M1r = 2'b00;
			14'b11110010000010: M1r = 2'b00;
			14'b00000110000010: M1r = 2'b01;
			14'b01000110000010: M1r = 2'b01;
			14'b10000110000010: M1r = 2'b10;
			14'b11000110000010: M1r = 2'b10;
			14'b00010110000010: M1r = 2'b01;
			14'b01010110000010: M1r = 2'b01;
			14'b10010110000010: M1r = 2'b01;
			14'b11010110000010: M1r = 2'b01;
			14'b00100110000010: M1r = 2'b00;
			14'b01100110000010: M1r = 2'b00;
			14'b10100110000010: M1r = 2'b01;
			14'b11100110000010: M1r = 2'b01;
			14'b00110110000010: M1r = 2'b00;
			14'b01110110000010: M1r = 2'b00;
			14'b10110110000010: M1r = 2'b00;
			14'b11110110000010: M1r = 2'b00;
			14'b00001010000010: M1r = 2'b10;
			14'b01001010000010: M1r = 2'b10;
			14'b10001010000010: M1r = 2'b10;
			14'b11001010000010: M1r = 2'b10;
			14'b00011010000010: M1r = 2'b10;
			14'b01011010000010: M1r = 2'b10;
			14'b10011010000010: M1r = 2'b10;
			14'b11011010000010: M1r = 2'b10;
			14'b00101010000010: M1r = 2'b01;
			14'b01101010000010: M1r = 2'b01;
			14'b10101010000010: M1r = 2'b01;
			14'b11101010000010: M1r = 2'b10;
			14'b00111010000010: M1r = 2'b01;
			14'b01111010000010: M1r = 2'b01;
			14'b10111010000010: M1r = 2'b01;
			14'b11111010000010: M1r = 2'b01;
			14'b00001110000010: M1r = 2'b11;
			14'b01001110000010: M1r = 2'b11;
			14'b10001110000010: M1r = 2'b11;
			14'b11001110000010: M1r = 2'b11;
			14'b00011110000010: M1r = 2'b10;
			14'b01011110000010: M1r = 2'b10;
			14'b10011110000010: M1r = 2'b11;
			14'b11011110000010: M1r = 2'b11;
			14'b00101110000010: M1r = 2'b10;
			14'b01101110000010: M1r = 2'b10;
			14'b10101110000010: M1r = 2'b10;
			14'b11101110000010: M1r = 2'b10;
			14'b00111110000010: M1r = 2'b01;
			14'b01111110000010: M1r = 2'b10;
			14'b10111110000010: M1r = 2'b10;
			14'b11111110000010: M1r = 2'b10;
			14'b00000011000010: M1r = 2'b00;
			14'b01000011000010: M1r = 2'b00;
			14'b10000011000010: M1r = 2'b01;
			14'b11000011000010: M1r = 2'b01;
			14'b00010011000010: M1r = 2'b00;
			14'b01010011000010: M1r = 2'b00;
			14'b10010011000010: M1r = 2'b00;
			14'b11010011000010: M1r = 2'b00;
			14'b00100011000010: M1r = 2'b00;
			14'b01100011000010: M1r = 2'b00;
			14'b10100011000010: M1r = 2'b00;
			14'b11100011000010: M1r = 2'b00;
			14'b00110011000010: M1r = 2'b00;
			14'b01110011000010: M1r = 2'b00;
			14'b10110011000010: M1r = 2'b00;
			14'b11110011000010: M1r = 2'b00;
			14'b00000111000010: M1r = 2'b01;
			14'b01000111000010: M1r = 2'b01;
			14'b10000111000010: M1r = 2'b01;
			14'b11000111000010: M1r = 2'b01;
			14'b00010111000010: M1r = 2'b01;
			14'b01010111000010: M1r = 2'b01;
			14'b10010111000010: M1r = 2'b01;
			14'b11010111000010: M1r = 2'b01;
			14'b00100111000010: M1r = 2'b00;
			14'b01100111000010: M1r = 2'b00;
			14'b10100111000010: M1r = 2'b00;
			14'b11100111000010: M1r = 2'b01;
			14'b00110111000010: M1r = 2'b00;
			14'b01110111000010: M1r = 2'b00;
			14'b10110111000010: M1r = 2'b00;
			14'b11110111000010: M1r = 2'b00;
			14'b00001011000010: M1r = 2'b10;
			14'b01001011000010: M1r = 2'b10;
			14'b10001011000010: M1r = 2'b10;
			14'b11001011000010: M1r = 2'b10;
			14'b00011011000010: M1r = 2'b01;
			14'b01011011000010: M1r = 2'b01;
			14'b10011011000010: M1r = 2'b10;
			14'b11011011000010: M1r = 2'b10;
			14'b00101011000010: M1r = 2'b01;
			14'b01101011000010: M1r = 2'b01;
			14'b10101011000010: M1r = 2'b01;
			14'b11101011000010: M1r = 2'b01;
			14'b00111011000010: M1r = 2'b00;
			14'b01111011000010: M1r = 2'b00;
			14'b10111011000010: M1r = 2'b01;
			14'b11111011000010: M1r = 2'b01;
			14'b00001111000010: M1r = 2'b10;
			14'b01001111000010: M1r = 2'b11;
			14'b10001111000010: M1r = 2'b11;
			14'b11001111000010: M1r = 2'b11;
			14'b00011111000010: M1r = 2'b10;
			14'b01011111000010: M1r = 2'b10;
			14'b10011111000010: M1r = 2'b10;
			14'b11011111000010: M1r = 2'b10;
			14'b00101111000010: M1r = 2'b10;
			14'b01101111000010: M1r = 2'b10;
			14'b10101111000010: M1r = 2'b10;
			14'b11101111000010: M1r = 2'b10;
			14'b00111111000010: M1r = 2'b01;
			14'b01111111000010: M1r = 2'b01;
			14'b10111111000010: M1r = 2'b01;
			14'b11111111000010: M1r = 2'b10;
			14'b00000000010010: M1r = 2'b10;
			14'b01000000010010: M1r = 2'b10;
			14'b10000000010010: M1r = 2'b10;
			14'b11000000010010: M1r = 2'b10;
			14'b00010000010010: M1r = 2'b01;
			14'b01010000010010: M1r = 2'b01;
			14'b10010000010010: M1r = 2'b01;
			14'b11010000010010: M1r = 2'b01;
			14'b00100000010010: M1r = 2'b01;
			14'b01100000010010: M1r = 2'b01;
			14'b10100000010010: M1r = 2'b01;
			14'b11100000010010: M1r = 2'b01;
			14'b00110000010010: M1r = 2'b00;
			14'b01110000010010: M1r = 2'b00;
			14'b10110000010010: M1r = 2'b00;
			14'b11110000010010: M1r = 2'b01;
			14'b00000100010010: M1r = 2'b10;
			14'b01000100010010: M1r = 2'b10;
			14'b10000100010010: M1r = 2'b11;
			14'b11000100010010: M1r = 2'b11;
			14'b00010100010010: M1r = 2'b10;
			14'b01010100010010: M1r = 2'b10;
			14'b10010100010010: M1r = 2'b10;
			14'b11010100010010: M1r = 2'b10;
			14'b00100100010010: M1r = 2'b01;
			14'b01100100010010: M1r = 2'b01;
			14'b10100100010010: M1r = 2'b10;
			14'b11100100010010: M1r = 2'b10;
			14'b00110100010010: M1r = 2'b01;
			14'b01110100010010: M1r = 2'b01;
			14'b10110100010010: M1r = 2'b01;
			14'b11110100010010: M1r = 2'b01;
			14'b00001000010010: M1r = 2'b11;
			14'b01001000010010: M1r = 2'b11;
			14'b10001000010010: M1r = 2'b11;
			14'b11001000010010: M1r = 2'b11;
			14'b00011000010010: M1r = 2'b11;
			14'b01011000010010: M1r = 2'b11;
			14'b10011000010010: M1r = 2'b11;
			14'b11011000010010: M1r = 2'b11;
			14'b00101000010010: M1r = 2'b10;
			14'b01101000010010: M1r = 2'b10;
			14'b10101000010010: M1r = 2'b10;
			14'b11101000010010: M1r = 2'b11;
			14'b00111000010010: M1r = 2'b10;
			14'b01111000010010: M1r = 2'b10;
			14'b10111000010010: M1r = 2'b10;
			14'b11111000010010: M1r = 2'b10;
			14'b00001100010010: M1r = 2'b11;
			14'b01001100010010: M1r = 2'b11;
			14'b10001100010010: M1r = 2'b11;
			14'b11001100010010: M1r = 2'b11;
			14'b00011100010010: M1r = 2'b11;
			14'b01011100010010: M1r = 2'b11;
			14'b10011100010010: M1r = 2'b11;
			14'b11011100010010: M1r = 2'b11;
			14'b00101100010010: M1r = 2'b11;
			14'b01101100010010: M1r = 2'b11;
			14'b10101100010010: M1r = 2'b11;
			14'b11101100010010: M1r = 2'b11;
			14'b00111100010010: M1r = 2'b10;
			14'b01111100010010: M1r = 2'b10;
			14'b10111100010010: M1r = 2'b11;
			14'b11111100010010: M1r = 2'b11;
			14'b00000001010010: M1r = 2'b01;
			14'b01000001010010: M1r = 2'b01;
			14'b10000001010010: M1r = 2'b10;
			14'b11000001010010: M1r = 2'b10;
			14'b00010001010010: M1r = 2'b01;
			14'b01010001010010: M1r = 2'b01;
			14'b10010001010010: M1r = 2'b01;
			14'b11010001010010: M1r = 2'b01;
			14'b00100001010010: M1r = 2'b00;
			14'b01100001010010: M1r = 2'b00;
			14'b10100001010010: M1r = 2'b01;
			14'b11100001010010: M1r = 2'b01;
			14'b00110001010010: M1r = 2'b00;
			14'b01110001010010: M1r = 2'b00;
			14'b10110001010010: M1r = 2'b00;
			14'b11110001010010: M1r = 2'b00;
			14'b00000101010010: M1r = 2'b10;
			14'b01000101010010: M1r = 2'b10;
			14'b10000101010010: M1r = 2'b10;
			14'b11000101010010: M1r = 2'b10;
			14'b00010101010010: M1r = 2'b10;
			14'b01010101010010: M1r = 2'b10;
			14'b10010101010010: M1r = 2'b10;
			14'b11010101010010: M1r = 2'b10;
			14'b00100101010010: M1r = 2'b01;
			14'b01100101010010: M1r = 2'b01;
			14'b10100101010010: M1r = 2'b01;
			14'b11100101010010: M1r = 2'b01;
			14'b00110101010010: M1r = 2'b01;
			14'b01110101010010: M1r = 2'b01;
			14'b10110101010010: M1r = 2'b01;
			14'b11110101010010: M1r = 2'b01;
			14'b00001001010010: M1r = 2'b11;
			14'b01001001010010: M1r = 2'b11;
			14'b10001001010010: M1r = 2'b11;
			14'b11001001010010: M1r = 2'b11;
			14'b00011001010010: M1r = 2'b10;
			14'b01011001010010: M1r = 2'b10;
			14'b10011001010010: M1r = 2'b11;
			14'b11011001010010: M1r = 2'b11;
			14'b00101001010010: M1r = 2'b10;
			14'b01101001010010: M1r = 2'b10;
			14'b10101001010010: M1r = 2'b10;
			14'b11101001010010: M1r = 2'b10;
			14'b00111001010010: M1r = 2'b01;
			14'b01111001010010: M1r = 2'b01;
			14'b10111001010010: M1r = 2'b10;
			14'b11111001010010: M1r = 2'b10;
			14'b00001101010010: M1r = 2'b11;
			14'b01001101010010: M1r = 2'b11;
			14'b10001101010010: M1r = 2'b11;
			14'b11001101010010: M1r = 2'b11;
			14'b00011101010010: M1r = 2'b11;
			14'b01011101010010: M1r = 2'b11;
			14'b10011101010010: M1r = 2'b11;
			14'b11011101010010: M1r = 2'b11;
			14'b00101101010010: M1r = 2'b11;
			14'b01101101010010: M1r = 2'b11;
			14'b10101101010010: M1r = 2'b11;
			14'b11101101010010: M1r = 2'b11;
			14'b00111101010010: M1r = 2'b10;
			14'b01111101010010: M1r = 2'b10;
			14'b10111101010010: M1r = 2'b10;
			14'b11111101010010: M1r = 2'b11;
			14'b00000010010010: M1r = 2'b01;
			14'b01000010010010: M1r = 2'b01;
			14'b10000010010010: M1r = 2'b01;
			14'b11000010010010: M1r = 2'b01;
			14'b00010010010010: M1r = 2'b00;
			14'b01010010010010: M1r = 2'b01;
			14'b10010010010010: M1r = 2'b01;
			14'b11010010010010: M1r = 2'b01;
			14'b00100010010010: M1r = 2'b00;
			14'b01100010010010: M1r = 2'b00;
			14'b10100010010010: M1r = 2'b00;
			14'b11100010010010: M1r = 2'b00;
			14'b00110010010010: M1r = 2'b00;
			14'b01110010010010: M1r = 2'b00;
			14'b10110010010010: M1r = 2'b00;
			14'b11110010010010: M1r = 2'b00;
			14'b00000110010010: M1r = 2'b10;
			14'b01000110010010: M1r = 2'b10;
			14'b10000110010010: M1r = 2'b10;
			14'b11000110010010: M1r = 2'b10;
			14'b00010110010010: M1r = 2'b01;
			14'b01010110010010: M1r = 2'b01;
			14'b10010110010010: M1r = 2'b10;
			14'b11010110010010: M1r = 2'b10;
			14'b00100110010010: M1r = 2'b01;
			14'b01100110010010: M1r = 2'b01;
			14'b10100110010010: M1r = 2'b01;
			14'b11100110010010: M1r = 2'b01;
			14'b00110110010010: M1r = 2'b00;
			14'b01110110010010: M1r = 2'b00;
			14'b10110110010010: M1r = 2'b01;
			14'b11110110010010: M1r = 2'b01;
			14'b00001010010010: M1r = 2'b10;
			14'b01001010010010: M1r = 2'b11;
			14'b10001010010010: M1r = 2'b11;
			14'b11001010010010: M1r = 2'b11;
			14'b00011010010010: M1r = 2'b10;
			14'b01011010010010: M1r = 2'b10;
			14'b10011010010010: M1r = 2'b10;
			14'b11011010010010: M1r = 2'b10;
			14'b00101010010010: M1r = 2'b10;
			14'b01101010010010: M1r = 2'b10;
			14'b10101010010010: M1r = 2'b10;
			14'b11101010010010: M1r = 2'b10;
			14'b00111010010010: M1r = 2'b01;
			14'b01111010010010: M1r = 2'b01;
			14'b10111010010010: M1r = 2'b01;
			14'b11111010010010: M1r = 2'b01;
			14'b00001110010010: M1r = 2'b11;
			14'b01001110010010: M1r = 2'b11;
			14'b10001110010010: M1r = 2'b11;
			14'b11001110010010: M1r = 2'b11;
			14'b00011110010010: M1r = 2'b11;
			14'b01011110010010: M1r = 2'b11;
			14'b10011110010010: M1r = 2'b11;
			14'b11011110010010: M1r = 2'b11;
			14'b00101110010010: M1r = 2'b10;
			14'b01101110010010: M1r = 2'b10;
			14'b10101110010010: M1r = 2'b11;
			14'b11101110010010: M1r = 2'b11;
			14'b00111110010010: M1r = 2'b10;
			14'b01111110010010: M1r = 2'b10;
			14'b10111110010010: M1r = 2'b10;
			14'b11111110010010: M1r = 2'b10;
			14'b00000011010010: M1r = 2'b01;
			14'b01000011010010: M1r = 2'b01;
			14'b10000011010010: M1r = 2'b01;
			14'b11000011010010: M1r = 2'b01;
			14'b00010011010010: M1r = 2'b00;
			14'b01010011010010: M1r = 2'b00;
			14'b10010011010010: M1r = 2'b01;
			14'b11010011010010: M1r = 2'b01;
			14'b00100011010010: M1r = 2'b00;
			14'b01100011010010: M1r = 2'b00;
			14'b10100011010010: M1r = 2'b00;
			14'b11100011010010: M1r = 2'b00;
			14'b00110011010010: M1r = 2'b00;
			14'b01110011010010: M1r = 2'b00;
			14'b10110011010010: M1r = 2'b00;
			14'b11110011010010: M1r = 2'b00;
			14'b00000111010010: M1r = 2'b01;
			14'b01000111010010: M1r = 2'b10;
			14'b10000111010010: M1r = 2'b10;
			14'b11000111010010: M1r = 2'b10;
			14'b00010111010010: M1r = 2'b01;
			14'b01010111010010: M1r = 2'b01;
			14'b10010111010010: M1r = 2'b01;
			14'b11010111010010: M1r = 2'b01;
			14'b00100111010010: M1r = 2'b00;
			14'b01100111010010: M1r = 2'b01;
			14'b10100111010010: M1r = 2'b01;
			14'b11100111010010: M1r = 2'b01;
			14'b00110111010010: M1r = 2'b00;
			14'b01110111010010: M1r = 2'b00;
			14'b10110111010010: M1r = 2'b00;
			14'b11110111010010: M1r = 2'b00;
			14'b00001011010010: M1r = 2'b10;
			14'b01001011010010: M1r = 2'b10;
			14'b10001011010010: M1r = 2'b10;
			14'b11001011010010: M1r = 2'b11;
			14'b00011011010010: M1r = 2'b10;
			14'b01011011010010: M1r = 2'b10;
			14'b10011011010010: M1r = 2'b10;
			14'b11011011010010: M1r = 2'b10;
			14'b00101011010010: M1r = 2'b01;
			14'b01101011010010: M1r = 2'b01;
			14'b10101011010010: M1r = 2'b10;
			14'b11101011010010: M1r = 2'b10;
			14'b00111011010010: M1r = 2'b01;
			14'b01111011010010: M1r = 2'b01;
			14'b10111011010010: M1r = 2'b01;
			14'b11111011010010: M1r = 2'b01;
			14'b00001111010010: M1r = 2'b11;
			14'b01001111010010: M1r = 2'b11;
			14'b10001111010010: M1r = 2'b11;
			14'b11001111010010: M1r = 2'b11;
			14'b00011111010010: M1r = 2'b10;
			14'b01011111010010: M1r = 2'b11;
			14'b10011111010010: M1r = 2'b11;
			14'b11011111010010: M1r = 2'b11;
			14'b00101111010010: M1r = 2'b10;
			14'b01101111010010: M1r = 2'b10;
			14'b10101111010010: M1r = 2'b10;
			14'b11101111010010: M1r = 2'b10;
			14'b00111111010010: M1r = 2'b10;
			14'b01111111010010: M1r = 2'b10;
			14'b10111111010010: M1r = 2'b10;
			14'b11111111010010: M1r = 2'b10;
			14'b00000000100010: M1r = 2'b10;
			14'b01000000100010: M1r = 2'b10;
			14'b10000000100010: M1r = 2'b10;
			14'b11000000100010: M1r = 2'b10;
			14'b00010000100010: M1r = 2'b01;
			14'b01010000100010: M1r = 2'b10;
			14'b10010000100010: M1r = 2'b10;
			14'b11010000100010: M1r = 2'b10;
			14'b00100000100010: M1r = 2'b01;
			14'b01100000100010: M1r = 2'b01;
			14'b10100000100010: M1r = 2'b01;
			14'b11100000100010: M1r = 2'b01;
			14'b00110000100010: M1r = 2'b01;
			14'b01110000100010: M1r = 2'b01;
			14'b10110000100010: M1r = 2'b01;
			14'b11110000100010: M1r = 2'b01;
			14'b00000100100010: M1r = 2'b11;
			14'b01000100100010: M1r = 2'b11;
			14'b10000100100010: M1r = 2'b11;
			14'b11000100100010: M1r = 2'b11;
			14'b00010100100010: M1r = 2'b10;
			14'b01010100100010: M1r = 2'b10;
			14'b10010100100010: M1r = 2'b11;
			14'b11010100100010: M1r = 2'b11;
			14'b00100100100010: M1r = 2'b10;
			14'b01100100100010: M1r = 2'b10;
			14'b10100100100010: M1r = 2'b10;
			14'b11100100100010: M1r = 2'b10;
			14'b00110100100010: M1r = 2'b01;
			14'b01110100100010: M1r = 2'b01;
			14'b10110100100010: M1r = 2'b10;
			14'b11110100100010: M1r = 2'b10;
			14'b00001000100010: M1r = 2'b11;
			14'b01001000100010: M1r = 2'b11;
			14'b10001000100010: M1r = 2'b11;
			14'b11001000100010: M1r = 2'b11;
			14'b00011000100010: M1r = 2'b11;
			14'b01011000100010: M1r = 2'b11;
			14'b10011000100010: M1r = 2'b11;
			14'b11011000100010: M1r = 2'b11;
			14'b00101000100010: M1r = 2'b10;
			14'b01101000100010: M1r = 2'b11;
			14'b10101000100010: M1r = 2'b11;
			14'b11101000100010: M1r = 2'b11;
			14'b00111000100010: M1r = 2'b10;
			14'b01111000100010: M1r = 2'b10;
			14'b10111000100010: M1r = 2'b10;
			14'b11111000100010: M1r = 2'b10;
			14'b00001100100010: M1r = 2'b11;
			14'b01001100100010: M1r = 2'b11;
			14'b10001100100010: M1r = 2'b11;
			14'b11001100100010: M1r = 2'b11;
			14'b00011100100010: M1r = 2'b11;
			14'b01011100100010: M1r = 2'b11;
			14'b10011100100010: M1r = 2'b11;
			14'b11011100100010: M1r = 2'b11;
			14'b00101100100010: M1r = 2'b11;
			14'b01101100100010: M1r = 2'b11;
			14'b10101100100010: M1r = 2'b11;
			14'b11101100100010: M1r = 2'b11;
			14'b00111100100010: M1r = 2'b11;
			14'b01111100100010: M1r = 2'b11;
			14'b10111100100010: M1r = 2'b11;
			14'b11111100100010: M1r = 2'b11;
			14'b00000001100010: M1r = 2'b10;
			14'b01000001100010: M1r = 2'b10;
			14'b10000001100010: M1r = 2'b10;
			14'b11000001100010: M1r = 2'b10;
			14'b00010001100010: M1r = 2'b01;
			14'b01010001100010: M1r = 2'b01;
			14'b10010001100010: M1r = 2'b01;
			14'b11010001100010: M1r = 2'b10;
			14'b00100001100010: M1r = 2'b01;
			14'b01100001100010: M1r = 2'b01;
			14'b10100001100010: M1r = 2'b01;
			14'b11100001100010: M1r = 2'b01;
			14'b00110001100010: M1r = 2'b00;
			14'b01110001100010: M1r = 2'b00;
			14'b10110001100010: M1r = 2'b01;
			14'b11110001100010: M1r = 2'b01;
			14'b00000101100010: M1r = 2'b10;
			14'b01000101100010: M1r = 2'b11;
			14'b10000101100010: M1r = 2'b11;
			14'b11000101100010: M1r = 2'b11;
			14'b00010101100010: M1r = 2'b10;
			14'b01010101100010: M1r = 2'b10;
			14'b10010101100010: M1r = 2'b10;
			14'b11010101100010: M1r = 2'b10;
			14'b00100101100010: M1r = 2'b01;
			14'b01100101100010: M1r = 2'b10;
			14'b10100101100010: M1r = 2'b10;
			14'b11100101100010: M1r = 2'b10;
			14'b00110101100010: M1r = 2'b01;
			14'b01110101100010: M1r = 2'b01;
			14'b10110101100010: M1r = 2'b01;
			14'b11110101100010: M1r = 2'b01;
			14'b00001001100010: M1r = 2'b11;
			14'b01001001100010: M1r = 2'b11;
			14'b10001001100010: M1r = 2'b11;
			14'b11001001100010: M1r = 2'b11;
			14'b00011001100010: M1r = 2'b11;
			14'b01011001100010: M1r = 2'b11;
			14'b10011001100010: M1r = 2'b11;
			14'b11011001100010: M1r = 2'b11;
			14'b00101001100010: M1r = 2'b10;
			14'b01101001100010: M1r = 2'b10;
			14'b10101001100010: M1r = 2'b11;
			14'b11101001100010: M1r = 2'b11;
			14'b00111001100010: M1r = 2'b10;
			14'b01111001100010: M1r = 2'b10;
			14'b10111001100010: M1r = 2'b10;
			14'b11111001100010: M1r = 2'b10;
			14'b00001101100010: M1r = 2'b11;
			14'b01001101100010: M1r = 2'b11;
			14'b10001101100010: M1r = 2'b11;
			14'b11001101100010: M1r = 2'b11;
			14'b00011101100010: M1r = 2'b11;
			14'b01011101100010: M1r = 2'b11;
			14'b10011101100010: M1r = 2'b11;
			14'b11011101100010: M1r = 2'b11;
			14'b00101101100010: M1r = 2'b11;
			14'b01101101100010: M1r = 2'b11;
			14'b10101101100010: M1r = 2'b11;
			14'b11101101100010: M1r = 2'b11;
			14'b00111101100010: M1r = 2'b10;
			14'b01111101100010: M1r = 2'b11;
			14'b10111101100010: M1r = 2'b11;
			14'b11111101100010: M1r = 2'b11;
			14'b00000010100010: M1r = 2'b01;
			14'b01000010100010: M1r = 2'b10;
			14'b10000010100010: M1r = 2'b10;
			14'b11000010100010: M1r = 2'b10;
			14'b00010010100010: M1r = 2'b01;
			14'b01010010100010: M1r = 2'b01;
			14'b10010010100010: M1r = 2'b01;
			14'b11010010100010: M1r = 2'b01;
			14'b00100010100010: M1r = 2'b00;
			14'b01100010100010: M1r = 2'b01;
			14'b10100010100010: M1r = 2'b01;
			14'b11100010100010: M1r = 2'b01;
			14'b00110010100010: M1r = 2'b00;
			14'b01110010100010: M1r = 2'b00;
			14'b10110010100010: M1r = 2'b00;
			14'b11110010100010: M1r = 2'b00;
			14'b00000110100010: M1r = 2'b10;
			14'b01000110100010: M1r = 2'b10;
			14'b10000110100010: M1r = 2'b10;
			14'b11000110100010: M1r = 2'b11;
			14'b00010110100010: M1r = 2'b10;
			14'b01010110100010: M1r = 2'b10;
			14'b10010110100010: M1r = 2'b10;
			14'b11010110100010: M1r = 2'b10;
			14'b00100110100010: M1r = 2'b01;
			14'b01100110100010: M1r = 2'b01;
			14'b10100110100010: M1r = 2'b01;
			14'b11100110100010: M1r = 2'b10;
			14'b00110110100010: M1r = 2'b01;
			14'b01110110100010: M1r = 2'b01;
			14'b10110110100010: M1r = 2'b01;
			14'b11110110100010: M1r = 2'b01;
			14'b00001010100010: M1r = 2'b11;
			14'b01001010100010: M1r = 2'b11;
			14'b10001010100010: M1r = 2'b11;
			14'b11001010100010: M1r = 2'b11;
			14'b00011010100010: M1r = 2'b10;
			14'b01011010100010: M1r = 2'b11;
			14'b10011010100010: M1r = 2'b11;
			14'b11011010100010: M1r = 2'b11;
			14'b00101010100010: M1r = 2'b10;
			14'b01101010100010: M1r = 2'b10;
			14'b10101010100010: M1r = 2'b10;
			14'b11101010100010: M1r = 2'b10;
			14'b00111010100010: M1r = 2'b01;
			14'b01111010100010: M1r = 2'b10;
			14'b10111010100010: M1r = 2'b10;
			14'b11111010100010: M1r = 2'b10;
			14'b00001110100010: M1r = 2'b11;
			14'b01001110100010: M1r = 2'b11;
			14'b10001110100010: M1r = 2'b11;
			14'b11001110100010: M1r = 2'b11;
			14'b00011110100010: M1r = 2'b11;
			14'b01011110100010: M1r = 2'b11;
			14'b10011110100010: M1r = 2'b11;
			14'b11011110100010: M1r = 2'b11;
			14'b00101110100010: M1r = 2'b11;
			14'b01101110100010: M1r = 2'b11;
			14'b10101110100010: M1r = 2'b11;
			14'b11101110100010: M1r = 2'b11;
			14'b00111110100010: M1r = 2'b10;
			14'b01111110100010: M1r = 2'b10;
			14'b10111110100010: M1r = 2'b11;
			14'b11111110100010: M1r = 2'b11;
			14'b00000011100010: M1r = 2'b01;
			14'b01000011100010: M1r = 2'b01;
			14'b10000011100010: M1r = 2'b01;
			14'b11000011100010: M1r = 2'b10;
			14'b00010011100010: M1r = 2'b01;
			14'b01010011100010: M1r = 2'b01;
			14'b10010011100010: M1r = 2'b01;
			14'b11010011100010: M1r = 2'b01;
			14'b00100011100010: M1r = 2'b00;
			14'b01100011100010: M1r = 2'b00;
			14'b10100011100010: M1r = 2'b00;
			14'b11100011100010: M1r = 2'b01;
			14'b00110011100010: M1r = 2'b00;
			14'b01110011100010: M1r = 2'b00;
			14'b10110011100010: M1r = 2'b00;
			14'b11110011100010: M1r = 2'b00;
			14'b00000111100010: M1r = 2'b10;
			14'b01000111100010: M1r = 2'b10;
			14'b10000111100010: M1r = 2'b10;
			14'b11000111100010: M1r = 2'b10;
			14'b00010111100010: M1r = 2'b01;
			14'b01010111100010: M1r = 2'b10;
			14'b10010111100010: M1r = 2'b10;
			14'b11010111100010: M1r = 2'b10;
			14'b00100111100010: M1r = 2'b01;
			14'b01100111100010: M1r = 2'b01;
			14'b10100111100010: M1r = 2'b01;
			14'b11100111100010: M1r = 2'b01;
			14'b00110111100010: M1r = 2'b00;
			14'b01110111100010: M1r = 2'b01;
			14'b10110111100010: M1r = 2'b01;
			14'b11110111100010: M1r = 2'b01;
			14'b00001011100010: M1r = 2'b11;
			14'b01001011100010: M1r = 2'b11;
			14'b10001011100010: M1r = 2'b11;
			14'b11001011100010: M1r = 2'b11;
			14'b00011011100010: M1r = 2'b10;
			14'b01011011100010: M1r = 2'b10;
			14'b10011011100010: M1r = 2'b10;
			14'b11011011100010: M1r = 2'b11;
			14'b00101011100010: M1r = 2'b10;
			14'b01101011100010: M1r = 2'b10;
			14'b10101011100010: M1r = 2'b10;
			14'b11101011100010: M1r = 2'b10;
			14'b00111011100010: M1r = 2'b01;
			14'b01111011100010: M1r = 2'b01;
			14'b10111011100010: M1r = 2'b01;
			14'b11111011100010: M1r = 2'b10;
			14'b00001111100010: M1r = 2'b11;
			14'b01001111100010: M1r = 2'b11;
			14'b10001111100010: M1r = 2'b11;
			14'b11001111100010: M1r = 2'b11;
			14'b00011111100010: M1r = 2'b11;
			14'b01011111100010: M1r = 2'b11;
			14'b10011111100010: M1r = 2'b11;
			14'b11011111100010: M1r = 2'b11;
			14'b00101111100010: M1r = 2'b10;
			14'b01101111100010: M1r = 2'b11;
			14'b10101111100010: M1r = 2'b11;
			14'b11101111100010: M1r = 2'b11;
			14'b00111111100010: M1r = 2'b10;
			14'b01111111100010: M1r = 2'b10;
			14'b10111111100010: M1r = 2'b10;
			14'b11111111100010: M1r = 2'b10;
			14'b00000000110010: M1r = 2'b10;
			14'b01000000110010: M1r = 2'b11;
			14'b10000000110010: M1r = 2'b11;
			14'b11000000110010: M1r = 2'b11;
			14'b00010000110010: M1r = 2'b10;
			14'b01010000110010: M1r = 2'b10;
			14'b10010000110010: M1r = 2'b10;
			14'b11010000110010: M1r = 2'b10;
			14'b00100000110010: M1r = 2'b01;
			14'b01100000110010: M1r = 2'b10;
			14'b10100000110010: M1r = 2'b10;
			14'b11100000110010: M1r = 2'b10;
			14'b00110000110010: M1r = 2'b01;
			14'b01110000110010: M1r = 2'b01;
			14'b10110000110010: M1r = 2'b01;
			14'b11110000110010: M1r = 2'b01;
			14'b00000100110010: M1r = 2'b11;
			14'b01000100110010: M1r = 2'b11;
			14'b10000100110010: M1r = 2'b11;
			14'b11000100110010: M1r = 2'b11;
			14'b00010100110010: M1r = 2'b11;
			14'b01010100110010: M1r = 2'b11;
			14'b10010100110010: M1r = 2'b11;
			14'b11010100110010: M1r = 2'b11;
			14'b00100100110010: M1r = 2'b10;
			14'b01100100110010: M1r = 2'b10;
			14'b10100100110010: M1r = 2'b10;
			14'b11100100110010: M1r = 2'b11;
			14'b00110100110010: M1r = 2'b10;
			14'b01110100110010: M1r = 2'b10;
			14'b10110100110010: M1r = 2'b10;
			14'b11110100110010: M1r = 2'b10;
			14'b00001000110010: M1r = 2'b11;
			14'b01001000110010: M1r = 2'b11;
			14'b10001000110010: M1r = 2'b11;
			14'b11001000110010: M1r = 2'b11;
			14'b00011000110010: M1r = 2'b11;
			14'b01011000110010: M1r = 2'b11;
			14'b10011000110010: M1r = 2'b11;
			14'b11011000110010: M1r = 2'b11;
			14'b00101000110010: M1r = 2'b11;
			14'b01101000110010: M1r = 2'b11;
			14'b10101000110010: M1r = 2'b11;
			14'b11101000110010: M1r = 2'b11;
			14'b00111000110010: M1r = 2'b10;
			14'b01111000110010: M1r = 2'b11;
			14'b10111000110010: M1r = 2'b11;
			14'b11111000110010: M1r = 2'b11;
			14'b00001100110010: M1r = 2'b11;
			14'b01001100110010: M1r = 2'b11;
			14'b10001100110010: M1r = 2'b11;
			14'b11001100110010: M1r = 2'b11;
			14'b00011100110010: M1r = 2'b11;
			14'b01011100110010: M1r = 2'b11;
			14'b10011100110010: M1r = 2'b11;
			14'b11011100110010: M1r = 2'b11;
			14'b00101100110010: M1r = 2'b11;
			14'b01101100110010: M1r = 2'b11;
			14'b10101100110010: M1r = 2'b11;
			14'b11101100110010: M1r = 2'b11;
			14'b00111100110010: M1r = 2'b11;
			14'b01111100110010: M1r = 2'b11;
			14'b10111100110010: M1r = 2'b11;
			14'b11111100110010: M1r = 2'b11;
			14'b00000001110010: M1r = 2'b10;
			14'b01000001110010: M1r = 2'b10;
			14'b10000001110010: M1r = 2'b10;
			14'b11000001110010: M1r = 2'b11;
			14'b00010001110010: M1r = 2'b10;
			14'b01010001110010: M1r = 2'b10;
			14'b10010001110010: M1r = 2'b10;
			14'b11010001110010: M1r = 2'b10;
			14'b00100001110010: M1r = 2'b01;
			14'b01100001110010: M1r = 2'b01;
			14'b10100001110010: M1r = 2'b01;
			14'b11100001110010: M1r = 2'b10;
			14'b00110001110010: M1r = 2'b01;
			14'b01110001110010: M1r = 2'b01;
			14'b10110001110010: M1r = 2'b01;
			14'b11110001110010: M1r = 2'b01;
			14'b00000101110010: M1r = 2'b11;
			14'b01000101110010: M1r = 2'b11;
			14'b10000101110010: M1r = 2'b11;
			14'b11000101110010: M1r = 2'b11;
			14'b00010101110010: M1r = 2'b10;
			14'b01010101110010: M1r = 2'b11;
			14'b10010101110010: M1r = 2'b11;
			14'b11010101110010: M1r = 2'b11;
			14'b00100101110010: M1r = 2'b10;
			14'b01100101110010: M1r = 2'b10;
			14'b10100101110010: M1r = 2'b10;
			14'b11100101110010: M1r = 2'b10;
			14'b00110101110010: M1r = 2'b01;
			14'b01110101110010: M1r = 2'b10;
			14'b10110101110010: M1r = 2'b10;
			14'b11110101110010: M1r = 2'b10;
			14'b00001001110010: M1r = 2'b11;
			14'b01001001110010: M1r = 2'b11;
			14'b10001001110010: M1r = 2'b11;
			14'b11001001110010: M1r = 2'b11;
			14'b00011001110010: M1r = 2'b11;
			14'b01011001110010: M1r = 2'b11;
			14'b10011001110010: M1r = 2'b11;
			14'b11011001110010: M1r = 2'b11;
			14'b00101001110010: M1r = 2'b11;
			14'b01101001110010: M1r = 2'b11;
			14'b10101001110010: M1r = 2'b11;
			14'b11101001110010: M1r = 2'b11;
			14'b00111001110010: M1r = 2'b10;
			14'b01111001110010: M1r = 2'b10;
			14'b10111001110010: M1r = 2'b10;
			14'b11111001110010: M1r = 2'b11;
			14'b00001101110010: M1r = 2'b11;
			14'b01001101110010: M1r = 2'b11;
			14'b10001101110010: M1r = 2'b11;
			14'b11001101110010: M1r = 2'b11;
			14'b00011101110010: M1r = 2'b11;
			14'b01011101110010: M1r = 2'b11;
			14'b10011101110010: M1r = 2'b11;
			14'b11011101110010: M1r = 2'b11;
			14'b00101101110010: M1r = 2'b11;
			14'b01101101110010: M1r = 2'b11;
			14'b10101101110010: M1r = 2'b11;
			14'b11101101110010: M1r = 2'b11;
			14'b00111101110010: M1r = 2'b11;
			14'b01111101110010: M1r = 2'b11;
			14'b10111101110010: M1r = 2'b11;
			14'b11111101110010: M1r = 2'b11;
			14'b00000010110010: M1r = 2'b10;
			14'b01000010110010: M1r = 2'b10;
			14'b10000010110010: M1r = 2'b10;
			14'b11000010110010: M1r = 2'b10;
			14'b00010010110010: M1r = 2'b01;
			14'b01010010110010: M1r = 2'b01;
			14'b10010010110010: M1r = 2'b10;
			14'b11010010110010: M1r = 2'b10;
			14'b00100010110010: M1r = 2'b01;
			14'b01100010110010: M1r = 2'b01;
			14'b10100010110010: M1r = 2'b01;
			14'b11100010110010: M1r = 2'b01;
			14'b00110010110010: M1r = 2'b00;
			14'b01110010110010: M1r = 2'b01;
			14'b10110010110010: M1r = 2'b01;
			14'b11110010110010: M1r = 2'b01;
			14'b00000110110010: M1r = 2'b11;
			14'b01000110110010: M1r = 2'b11;
			14'b10000110110010: M1r = 2'b11;
			14'b11000110110010: M1r = 2'b11;
			14'b00010110110010: M1r = 2'b10;
			14'b01010110110010: M1r = 2'b10;
			14'b10010110110010: M1r = 2'b10;
			14'b11010110110010: M1r = 2'b11;
			14'b00100110110010: M1r = 2'b10;
			14'b01100110110010: M1r = 2'b10;
			14'b10100110110010: M1r = 2'b10;
			14'b11100110110010: M1r = 2'b10;
			14'b00110110110010: M1r = 2'b01;
			14'b01110110110010: M1r = 2'b01;
			14'b10110110110010: M1r = 2'b01;
			14'b11110110110010: M1r = 2'b10;
			14'b00001010110010: M1r = 2'b11;
			14'b01001010110010: M1r = 2'b11;
			14'b10001010110010: M1r = 2'b11;
			14'b11001010110010: M1r = 2'b11;
			14'b00011010110010: M1r = 2'b11;
			14'b01011010110010: M1r = 2'b11;
			14'b10011010110010: M1r = 2'b11;
			14'b11011010110010: M1r = 2'b11;
			14'b00101010110010: M1r = 2'b10;
			14'b01101010110010: M1r = 2'b11;
			14'b10101010110010: M1r = 2'b11;
			14'b11101010110010: M1r = 2'b11;
			14'b00111010110010: M1r = 2'b10;
			14'b01111010110010: M1r = 2'b10;
			14'b10111010110010: M1r = 2'b10;
			14'b11111010110010: M1r = 2'b10;
			14'b00001110110010: M1r = 2'b11;
			14'b01001110110010: M1r = 2'b11;
			14'b10001110110010: M1r = 2'b11;
			14'b11001110110010: M1r = 2'b11;
			14'b00011110110010: M1r = 2'b11;
			14'b01011110110010: M1r = 2'b11;
			14'b10011110110010: M1r = 2'b11;
			14'b11011110110010: M1r = 2'b11;
			14'b00101110110010: M1r = 2'b11;
			14'b01101110110010: M1r = 2'b11;
			14'b10101110110010: M1r = 2'b11;
			14'b11101110110010: M1r = 2'b11;
			14'b00111110110010: M1r = 2'b11;
			14'b01111110110010: M1r = 2'b11;
			14'b10111110110010: M1r = 2'b11;
			14'b11111110110010: M1r = 2'b11;
			14'b00000011110010: M1r = 2'b10;
			14'b01000011110010: M1r = 2'b10;
			14'b10000011110010: M1r = 2'b10;
			14'b11000011110010: M1r = 2'b10;
			14'b00010011110010: M1r = 2'b01;
			14'b01010011110010: M1r = 2'b01;
			14'b10010011110010: M1r = 2'b01;
			14'b11010011110010: M1r = 2'b10;
			14'b00100011110010: M1r = 2'b01;
			14'b01100011110010: M1r = 2'b01;
			14'b10100011110010: M1r = 2'b01;
			14'b11100011110010: M1r = 2'b01;
			14'b00110011110010: M1r = 2'b00;
			14'b01110011110010: M1r = 2'b00;
			14'b10110011110010: M1r = 2'b00;
			14'b11110011110010: M1r = 2'b01;
			14'b00000111110010: M1r = 2'b10;
			14'b01000111110010: M1r = 2'b10;
			14'b10000111110010: M1r = 2'b11;
			14'b11000111110010: M1r = 2'b11;
			14'b00010111110010: M1r = 2'b10;
			14'b01010111110010: M1r = 2'b10;
			14'b10010111110010: M1r = 2'b10;
			14'b11010111110010: M1r = 2'b10;
			14'b00100111110010: M1r = 2'b01;
			14'b01100111110010: M1r = 2'b01;
			14'b10100111110010: M1r = 2'b10;
			14'b11100111110010: M1r = 2'b10;
			14'b00110111110010: M1r = 2'b01;
			14'b01110111110010: M1r = 2'b01;
			14'b10110111110010: M1r = 2'b01;
			14'b11110111110010: M1r = 2'b01;
			14'b00001011110010: M1r = 2'b11;
			14'b01001011110010: M1r = 2'b11;
			14'b10001011110010: M1r = 2'b11;
			14'b11001011110010: M1r = 2'b11;
			14'b00011011110010: M1r = 2'b11;
			14'b01011011110010: M1r = 2'b11;
			14'b10011011110010: M1r = 2'b11;
			14'b11011011110010: M1r = 2'b11;
			14'b00101011110010: M1r = 2'b10;
			14'b01101011110010: M1r = 2'b10;
			14'b10101011110010: M1r = 2'b10;
			14'b11101011110010: M1r = 2'b11;
			14'b00111011110010: M1r = 2'b10;
			14'b01111011110010: M1r = 2'b10;
			14'b10111011110010: M1r = 2'b10;
			14'b11111011110010: M1r = 2'b10;
			14'b00001111110010: M1r = 2'b11;
			14'b01001111110010: M1r = 2'b11;
			14'b10001111110010: M1r = 2'b11;
			14'b11001111110010: M1r = 2'b11;
			14'b00011111110010: M1r = 2'b11;
			14'b01011111110010: M1r = 2'b11;
			14'b10011111110010: M1r = 2'b11;
			14'b11011111110010: M1r = 2'b11;
			14'b00101111110010: M1r = 2'b11;
			14'b01101111110010: M1r = 2'b11;
			14'b10101111110010: M1r = 2'b11;
			14'b11101111110010: M1r = 2'b11;
			14'b00111111110010: M1r = 2'b10;
			14'b01111111110010: M1r = 2'b11;
			14'b10111111110010: M1r = 2'b11;
			14'b11111111110010: M1r = 2'b11;
			14'b00000000000110: M1r = 2'b00;
			14'b01000000000110: M1r = 2'b00;
			14'b10000000000110: M1r = 2'b01;
			14'b11000000000110: M1r = 2'b01;
			14'b00010000000110: M1r = 2'b00;
			14'b01010000000110: M1r = 2'b00;
			14'b10010000000110: M1r = 2'b00;
			14'b11010000000110: M1r = 2'b00;
			14'b00100000000110: M1r = 2'b00;
			14'b01100000000110: M1r = 2'b00;
			14'b10100000000110: M1r = 2'b00;
			14'b11100000000110: M1r = 2'b00;
			14'b00110000000110: M1r = 2'b00;
			14'b01110000000110: M1r = 2'b00;
			14'b10110000000110: M1r = 2'b00;
			14'b11110000000110: M1r = 2'b00;
			14'b00000100000110: M1r = 2'b01;
			14'b01000100000110: M1r = 2'b01;
			14'b10000100000110: M1r = 2'b01;
			14'b11000100000110: M1r = 2'b10;
			14'b00010100000110: M1r = 2'b01;
			14'b01010100000110: M1r = 2'b01;
			14'b10010100000110: M1r = 2'b01;
			14'b11010100000110: M1r = 2'b01;
			14'b00100100000110: M1r = 2'b00;
			14'b01100100000110: M1r = 2'b00;
			14'b10100100000110: M1r = 2'b00;
			14'b11100100000110: M1r = 2'b01;
			14'b00110100000110: M1r = 2'b00;
			14'b01110100000110: M1r = 2'b00;
			14'b10110100000110: M1r = 2'b00;
			14'b11110100000110: M1r = 2'b00;
			14'b00001000000110: M1r = 2'b10;
			14'b01001000000110: M1r = 2'b10;
			14'b10001000000110: M1r = 2'b10;
			14'b11001000000110: M1r = 2'b10;
			14'b00011000000110: M1r = 2'b01;
			14'b01011000000110: M1r = 2'b01;
			14'b10011000000110: M1r = 2'b10;
			14'b11011000000110: M1r = 2'b10;
			14'b00101000000110: M1r = 2'b01;
			14'b01101000000110: M1r = 2'b01;
			14'b10101000000110: M1r = 2'b01;
			14'b11101000000110: M1r = 2'b01;
			14'b00111000000110: M1r = 2'b00;
			14'b01111000000110: M1r = 2'b01;
			14'b10111000000110: M1r = 2'b01;
			14'b11111000000110: M1r = 2'b01;
			14'b00001100000110: M1r = 2'b11;
			14'b01001100000110: M1r = 2'b11;
			14'b10001100000110: M1r = 2'b11;
			14'b11001100000110: M1r = 2'b11;
			14'b00011100000110: M1r = 2'b10;
			14'b01011100000110: M1r = 2'b10;
			14'b10011100000110: M1r = 2'b10;
			14'b11011100000110: M1r = 2'b11;
			14'b00101100000110: M1r = 2'b10;
			14'b01101100000110: M1r = 2'b10;
			14'b10101100000110: M1r = 2'b10;
			14'b11101100000110: M1r = 2'b10;
			14'b00111100000110: M1r = 2'b01;
			14'b01111100000110: M1r = 2'b01;
			14'b10111100000110: M1r = 2'b01;
			14'b11111100000110: M1r = 2'b10;
			14'b00000001000110: M1r = 2'b00;
			14'b01000001000110: M1r = 2'b00;
			14'b10000001000110: M1r = 2'b00;
			14'b11000001000110: M1r = 2'b00;
			14'b00010001000110: M1r = 2'b00;
			14'b01010001000110: M1r = 2'b00;
			14'b10010001000110: M1r = 2'b00;
			14'b11010001000110: M1r = 2'b00;
			14'b00100001000110: M1r = 2'b00;
			14'b01100001000110: M1r = 2'b00;
			14'b10100001000110: M1r = 2'b00;
			14'b11100001000110: M1r = 2'b00;
			14'b00110001000110: M1r = 2'b00;
			14'b01110001000110: M1r = 2'b00;
			14'b10110001000110: M1r = 2'b00;
			14'b11110001000110: M1r = 2'b00;
			14'b00000101000110: M1r = 2'b01;
			14'b01000101000110: M1r = 2'b01;
			14'b10000101000110: M1r = 2'b01;
			14'b11000101000110: M1r = 2'b01;
			14'b00010101000110: M1r = 2'b00;
			14'b01010101000110: M1r = 2'b00;
			14'b10010101000110: M1r = 2'b01;
			14'b11010101000110: M1r = 2'b01;
			14'b00100101000110: M1r = 2'b00;
			14'b01100101000110: M1r = 2'b00;
			14'b10100101000110: M1r = 2'b00;
			14'b11100101000110: M1r = 2'b00;
			14'b00110101000110: M1r = 2'b00;
			14'b01110101000110: M1r = 2'b00;
			14'b10110101000110: M1r = 2'b00;
			14'b11110101000110: M1r = 2'b00;
			14'b00001001000110: M1r = 2'b10;
			14'b01001001000110: M1r = 2'b10;
			14'b10001001000110: M1r = 2'b10;
			14'b11001001000110: M1r = 2'b10;
			14'b00011001000110: M1r = 2'b01;
			14'b01011001000110: M1r = 2'b01;
			14'b10011001000110: M1r = 2'b01;
			14'b11011001000110: M1r = 2'b10;
			14'b00101001000110: M1r = 2'b01;
			14'b01101001000110: M1r = 2'b01;
			14'b10101001000110: M1r = 2'b01;
			14'b11101001000110: M1r = 2'b01;
			14'b00111001000110: M1r = 2'b00;
			14'b01111001000110: M1r = 2'b00;
			14'b10111001000110: M1r = 2'b00;
			14'b11111001000110: M1r = 2'b01;
			14'b00001101000110: M1r = 2'b10;
			14'b01001101000110: M1r = 2'b10;
			14'b10001101000110: M1r = 2'b11;
			14'b11001101000110: M1r = 2'b11;
			14'b00011101000110: M1r = 2'b10;
			14'b01011101000110: M1r = 2'b10;
			14'b10011101000110: M1r = 2'b10;
			14'b11011101000110: M1r = 2'b10;
			14'b00101101000110: M1r = 2'b01;
			14'b01101101000110: M1r = 2'b01;
			14'b10101101000110: M1r = 2'b10;
			14'b11101101000110: M1r = 2'b10;
			14'b00111101000110: M1r = 2'b01;
			14'b01111101000110: M1r = 2'b01;
			14'b10111101000110: M1r = 2'b01;
			14'b11111101000110: M1r = 2'b01;
			14'b00000010000110: M1r = 2'b00;
			14'b01000010000110: M1r = 2'b00;
			14'b10000010000110: M1r = 2'b00;
			14'b11000010000110: M1r = 2'b00;
			14'b00010010000110: M1r = 2'b00;
			14'b01010010000110: M1r = 2'b00;
			14'b10010010000110: M1r = 2'b00;
			14'b11010010000110: M1r = 2'b00;
			14'b00100010000110: M1r = 2'b00;
			14'b01100010000110: M1r = 2'b00;
			14'b10100010000110: M1r = 2'b00;
			14'b11100010000110: M1r = 2'b00;
			14'b00110010000110: M1r = 2'b00;
			14'b01110010000110: M1r = 2'b00;
			14'b10110010000110: M1r = 2'b00;
			14'b11110010000110: M1r = 2'b00;
			14'b00000110000110: M1r = 2'b00;
			14'b01000110000110: M1r = 2'b01;
			14'b10000110000110: M1r = 2'b01;
			14'b11000110000110: M1r = 2'b01;
			14'b00010110000110: M1r = 2'b00;
			14'b01010110000110: M1r = 2'b00;
			14'b10010110000110: M1r = 2'b00;
			14'b11010110000110: M1r = 2'b00;
			14'b00100110000110: M1r = 2'b00;
			14'b01100110000110: M1r = 2'b00;
			14'b10100110000110: M1r = 2'b00;
			14'b11100110000110: M1r = 2'b00;
			14'b00110110000110: M1r = 2'b00;
			14'b01110110000110: M1r = 2'b00;
			14'b10110110000110: M1r = 2'b00;
			14'b11110110000110: M1r = 2'b00;
			14'b00001010000110: M1r = 2'b01;
			14'b01001010000110: M1r = 2'b01;
			14'b10001010000110: M1r = 2'b10;
			14'b11001010000110: M1r = 2'b10;
			14'b00011010000110: M1r = 2'b01;
			14'b01011010000110: M1r = 2'b01;
			14'b10011010000110: M1r = 2'b01;
			14'b11011010000110: M1r = 2'b01;
			14'b00101010000110: M1r = 2'b00;
			14'b01101010000110: M1r = 2'b00;
			14'b10101010000110: M1r = 2'b01;
			14'b11101010000110: M1r = 2'b01;
			14'b00111010000110: M1r = 2'b00;
			14'b01111010000110: M1r = 2'b00;
			14'b10111010000110: M1r = 2'b00;
			14'b11111010000110: M1r = 2'b00;
			14'b00001110000110: M1r = 2'b10;
			14'b01001110000110: M1r = 2'b10;
			14'b10001110000110: M1r = 2'b10;
			14'b11001110000110: M1r = 2'b10;
			14'b00011110000110: M1r = 2'b10;
			14'b01011110000110: M1r = 2'b10;
			14'b10011110000110: M1r = 2'b10;
			14'b11011110000110: M1r = 2'b10;
			14'b00101110000110: M1r = 2'b01;
			14'b01101110000110: M1r = 2'b01;
			14'b10101110000110: M1r = 2'b01;
			14'b11101110000110: M1r = 2'b10;
			14'b00111110000110: M1r = 2'b01;
			14'b01111110000110: M1r = 2'b01;
			14'b10111110000110: M1r = 2'b01;
			14'b11111110000110: M1r = 2'b01;
			14'b00000011000110: M1r = 2'b00;
			14'b01000011000110: M1r = 2'b00;
			14'b10000011000110: M1r = 2'b00;
			14'b11000011000110: M1r = 2'b00;
			14'b00010011000110: M1r = 2'b00;
			14'b01010011000110: M1r = 2'b00;
			14'b10010011000110: M1r = 2'b00;
			14'b11010011000110: M1r = 2'b00;
			14'b00100011000110: M1r = 2'b00;
			14'b01100011000110: M1r = 2'b00;
			14'b10100011000110: M1r = 2'b00;
			14'b11100011000110: M1r = 2'b00;
			14'b00110011000110: M1r = 2'b00;
			14'b01110011000110: M1r = 2'b00;
			14'b10110011000110: M1r = 2'b00;
			14'b11110011000110: M1r = 2'b00;
			14'b00000111000110: M1r = 2'b00;
			14'b01000111000110: M1r = 2'b00;
			14'b10000111000110: M1r = 2'b01;
			14'b11000111000110: M1r = 2'b01;
			14'b00010111000110: M1r = 2'b00;
			14'b01010111000110: M1r = 2'b00;
			14'b10010111000110: M1r = 2'b00;
			14'b11010111000110: M1r = 2'b00;
			14'b00100111000110: M1r = 2'b00;
			14'b01100111000110: M1r = 2'b00;
			14'b10100111000110: M1r = 2'b00;
			14'b11100111000110: M1r = 2'b00;
			14'b00110111000110: M1r = 2'b00;
			14'b01110111000110: M1r = 2'b00;
			14'b10110111000110: M1r = 2'b00;
			14'b11110111000110: M1r = 2'b00;
			14'b00001011000110: M1r = 2'b01;
			14'b01001011000110: M1r = 2'b01;
			14'b10001011000110: M1r = 2'b01;
			14'b11001011000110: M1r = 2'b01;
			14'b00011011000110: M1r = 2'b00;
			14'b01011011000110: M1r = 2'b01;
			14'b10011011000110: M1r = 2'b01;
			14'b11011011000110: M1r = 2'b01;
			14'b00101011000110: M1r = 2'b00;
			14'b01101011000110: M1r = 2'b00;
			14'b10101011000110: M1r = 2'b00;
			14'b11101011000110: M1r = 2'b00;
			14'b00111011000110: M1r = 2'b00;
			14'b01111011000110: M1r = 2'b00;
			14'b10111011000110: M1r = 2'b00;
			14'b11111011000110: M1r = 2'b00;
			14'b00001111000110: M1r = 2'b10;
			14'b01001111000110: M1r = 2'b10;
			14'b10001111000110: M1r = 2'b10;
			14'b11001111000110: M1r = 2'b10;
			14'b00011111000110: M1r = 2'b01;
			14'b01011111000110: M1r = 2'b01;
			14'b10011111000110: M1r = 2'b10;
			14'b11011111000110: M1r = 2'b10;
			14'b00101111000110: M1r = 2'b01;
			14'b01101111000110: M1r = 2'b01;
			14'b10101111000110: M1r = 2'b01;
			14'b11101111000110: M1r = 2'b01;
			14'b00111111000110: M1r = 2'b00;
			14'b01111111000110: M1r = 2'b00;
			14'b10111111000110: M1r = 2'b01;
			14'b11111111000110: M1r = 2'b01;
			14'b00000000010110: M1r = 2'b01;
			14'b01000000010110: M1r = 2'b01;
			14'b10000000010110: M1r = 2'b01;
			14'b11000000010110: M1r = 2'b01;
			14'b00010000010110: M1r = 2'b00;
			14'b01010000010110: M1r = 2'b00;
			14'b10010000010110: M1r = 2'b01;
			14'b11010000010110: M1r = 2'b01;
			14'b00100000010110: M1r = 2'b00;
			14'b01100000010110: M1r = 2'b00;
			14'b10100000010110: M1r = 2'b00;
			14'b11100000010110: M1r = 2'b00;
			14'b00110000010110: M1r = 2'b00;
			14'b01110000010110: M1r = 2'b00;
			14'b10110000010110: M1r = 2'b00;
			14'b11110000010110: M1r = 2'b00;
			14'b00000100010110: M1r = 2'b01;
			14'b01000100010110: M1r = 2'b10;
			14'b10000100010110: M1r = 2'b10;
			14'b11000100010110: M1r = 2'b10;
			14'b00010100010110: M1r = 2'b01;
			14'b01010100010110: M1r = 2'b01;
			14'b10010100010110: M1r = 2'b01;
			14'b11010100010110: M1r = 2'b01;
			14'b00100100010110: M1r = 2'b01;
			14'b01100100010110: M1r = 2'b01;
			14'b10100100010110: M1r = 2'b01;
			14'b11100100010110: M1r = 2'b01;
			14'b00110100010110: M1r = 2'b00;
			14'b01110100010110: M1r = 2'b00;
			14'b10110100010110: M1r = 2'b00;
			14'b11110100010110: M1r = 2'b01;
			14'b00001000010110: M1r = 2'b10;
			14'b01001000010110: M1r = 2'b10;
			14'b10001000010110: M1r = 2'b11;
			14'b11001000010110: M1r = 2'b11;
			14'b00011000010110: M1r = 2'b10;
			14'b01011000010110: M1r = 2'b10;
			14'b10011000010110: M1r = 2'b10;
			14'b11011000010110: M1r = 2'b10;
			14'b00101000010110: M1r = 2'b01;
			14'b01101000010110: M1r = 2'b01;
			14'b10101000010110: M1r = 2'b10;
			14'b11101000010110: M1r = 2'b10;
			14'b00111000010110: M1r = 2'b01;
			14'b01111000010110: M1r = 2'b01;
			14'b10111000010110: M1r = 2'b01;
			14'b11111000010110: M1r = 2'b01;
			14'b00001100010110: M1r = 2'b11;
			14'b01001100010110: M1r = 2'b11;
			14'b10001100010110: M1r = 2'b11;
			14'b11001100010110: M1r = 2'b11;
			14'b00011100010110: M1r = 2'b11;
			14'b01011100010110: M1r = 2'b11;
			14'b10011100010110: M1r = 2'b11;
			14'b11011100010110: M1r = 2'b11;
			14'b00101100010110: M1r = 2'b10;
			14'b01101100010110: M1r = 2'b10;
			14'b10101100010110: M1r = 2'b10;
			14'b11101100010110: M1r = 2'b10;
			14'b00111100010110: M1r = 2'b10;
			14'b01111100010110: M1r = 2'b10;
			14'b10111100010110: M1r = 2'b10;
			14'b11111100010110: M1r = 2'b10;
			14'b00000001010110: M1r = 2'b00;
			14'b01000001010110: M1r = 2'b01;
			14'b10000001010110: M1r = 2'b01;
			14'b11000001010110: M1r = 2'b01;
			14'b00010001010110: M1r = 2'b00;
			14'b01010001010110: M1r = 2'b00;
			14'b10010001010110: M1r = 2'b00;
			14'b11010001010110: M1r = 2'b00;
			14'b00100001010110: M1r = 2'b00;
			14'b01100001010110: M1r = 2'b00;
			14'b10100001010110: M1r = 2'b00;
			14'b11100001010110: M1r = 2'b00;
			14'b00110001010110: M1r = 2'b00;
			14'b01110001010110: M1r = 2'b00;
			14'b10110001010110: M1r = 2'b00;
			14'b11110001010110: M1r = 2'b00;
			14'b00000101010110: M1r = 2'b01;
			14'b01000101010110: M1r = 2'b01;
			14'b10000101010110: M1r = 2'b10;
			14'b11000101010110: M1r = 2'b10;
			14'b00010101010110: M1r = 2'b01;
			14'b01010101010110: M1r = 2'b01;
			14'b10010101010110: M1r = 2'b01;
			14'b11010101010110: M1r = 2'b01;
			14'b00100101010110: M1r = 2'b00;
			14'b01100101010110: M1r = 2'b00;
			14'b10100101010110: M1r = 2'b01;
			14'b11100101010110: M1r = 2'b01;
			14'b00110101010110: M1r = 2'b00;
			14'b01110101010110: M1r = 2'b00;
			14'b10110101010110: M1r = 2'b00;
			14'b11110101010110: M1r = 2'b00;
			14'b00001001010110: M1r = 2'b10;
			14'b01001001010110: M1r = 2'b10;
			14'b10001001010110: M1r = 2'b10;
			14'b11001001010110: M1r = 2'b10;
			14'b00011001010110: M1r = 2'b01;
			14'b01011001010110: M1r = 2'b10;
			14'b10011001010110: M1r = 2'b10;
			14'b11011001010110: M1r = 2'b10;
			14'b00101001010110: M1r = 2'b01;
			14'b01101001010110: M1r = 2'b01;
			14'b10101001010110: M1r = 2'b01;
			14'b11101001010110: M1r = 2'b01;
			14'b00111001010110: M1r = 2'b01;
			14'b01111001010110: M1r = 2'b01;
			14'b10111001010110: M1r = 2'b01;
			14'b11111001010110: M1r = 2'b01;
			14'b00001101010110: M1r = 2'b11;
			14'b01001101010110: M1r = 2'b11;
			14'b10001101010110: M1r = 2'b11;
			14'b11001101010110: M1r = 2'b11;
			14'b00011101010110: M1r = 2'b10;
			14'b01011101010110: M1r = 2'b10;
			14'b10011101010110: M1r = 2'b11;
			14'b11011101010110: M1r = 2'b11;
			14'b00101101010110: M1r = 2'b10;
			14'b01101101010110: M1r = 2'b10;
			14'b10101101010110: M1r = 2'b10;
			14'b11101101010110: M1r = 2'b10;
			14'b00111101010110: M1r = 2'b01;
			14'b01111101010110: M1r = 2'b01;
			14'b10111101010110: M1r = 2'b10;
			14'b11111101010110: M1r = 2'b10;
			14'b00000010010110: M1r = 2'b00;
			14'b01000010010110: M1r = 2'b00;
			14'b10000010010110: M1r = 2'b00;
			14'b11000010010110: M1r = 2'b01;
			14'b00010010010110: M1r = 2'b00;
			14'b01010010010110: M1r = 2'b00;
			14'b10010010010110: M1r = 2'b00;
			14'b11010010010110: M1r = 2'b00;
			14'b00100010010110: M1r = 2'b00;
			14'b01100010010110: M1r = 2'b00;
			14'b10100010010110: M1r = 2'b00;
			14'b11100010010110: M1r = 2'b00;
			14'b00110010010110: M1r = 2'b00;
			14'b01110010010110: M1r = 2'b00;
			14'b10110010010110: M1r = 2'b00;
			14'b11110010010110: M1r = 2'b00;
			14'b00000110010110: M1r = 2'b01;
			14'b01000110010110: M1r = 2'b01;
			14'b10000110010110: M1r = 2'b01;
			14'b11000110010110: M1r = 2'b01;
			14'b00010110010110: M1r = 2'b00;
			14'b01010110010110: M1r = 2'b01;
			14'b10010110010110: M1r = 2'b01;
			14'b11010110010110: M1r = 2'b01;
			14'b00100110010110: M1r = 2'b00;
			14'b01100110010110: M1r = 2'b00;
			14'b10100110010110: M1r = 2'b00;
			14'b11100110010110: M1r = 2'b00;
			14'b00110110010110: M1r = 2'b00;
			14'b01110110010110: M1r = 2'b00;
			14'b10110110010110: M1r = 2'b00;
			14'b11110110010110: M1r = 2'b00;
			14'b00001010010110: M1r = 2'b10;
			14'b01001010010110: M1r = 2'b10;
			14'b10001010010110: M1r = 2'b10;
			14'b11001010010110: M1r = 2'b10;
			14'b00011010010110: M1r = 2'b01;
			14'b01011010010110: M1r = 2'b01;
			14'b10011010010110: M1r = 2'b10;
			14'b11011010010110: M1r = 2'b10;
			14'b00101010010110: M1r = 2'b01;
			14'b01101010010110: M1r = 2'b01;
			14'b10101010010110: M1r = 2'b01;
			14'b11101010010110: M1r = 2'b01;
			14'b00111010010110: M1r = 2'b00;
			14'b01111010010110: M1r = 2'b00;
			14'b10111010010110: M1r = 2'b01;
			14'b11111010010110: M1r = 2'b01;
			14'b00001110010110: M1r = 2'b10;
			14'b01001110010110: M1r = 2'b11;
			14'b10001110010110: M1r = 2'b11;
			14'b11001110010110: M1r = 2'b11;
			14'b00011110010110: M1r = 2'b10;
			14'b01011110010110: M1r = 2'b10;
			14'b10011110010110: M1r = 2'b10;
			14'b11011110010110: M1r = 2'b10;
			14'b00101110010110: M1r = 2'b01;
			14'b01101110010110: M1r = 2'b10;
			14'b10101110010110: M1r = 2'b10;
			14'b11101110010110: M1r = 2'b10;
			14'b00111110010110: M1r = 2'b01;
			14'b01111110010110: M1r = 2'b01;
			14'b10111110010110: M1r = 2'b01;
			14'b11111110010110: M1r = 2'b01;
			14'b00000011010110: M1r = 2'b00;
			14'b01000011010110: M1r = 2'b00;
			14'b10000011010110: M1r = 2'b00;
			14'b11000011010110: M1r = 2'b00;
			14'b00010011010110: M1r = 2'b00;
			14'b01010011010110: M1r = 2'b00;
			14'b10010011010110: M1r = 2'b00;
			14'b11010011010110: M1r = 2'b00;
			14'b00100011010110: M1r = 2'b00;
			14'b01100011010110: M1r = 2'b00;
			14'b10100011010110: M1r = 2'b00;
			14'b11100011010110: M1r = 2'b00;
			14'b00110011010110: M1r = 2'b00;
			14'b01110011010110: M1r = 2'b00;
			14'b10110011010110: M1r = 2'b00;
			14'b11110011010110: M1r = 2'b00;
			14'b00000111010110: M1r = 2'b01;
			14'b01000111010110: M1r = 2'b01;
			14'b10000111010110: M1r = 2'b01;
			14'b11000111010110: M1r = 2'b01;
			14'b00010111010110: M1r = 2'b00;
			14'b01010111010110: M1r = 2'b00;
			14'b10010111010110: M1r = 2'b00;
			14'b11010111010110: M1r = 2'b01;
			14'b00100111010110: M1r = 2'b00;
			14'b01100111010110: M1r = 2'b00;
			14'b10100111010110: M1r = 2'b00;
			14'b11100111010110: M1r = 2'b00;
			14'b00110111010110: M1r = 2'b00;
			14'b01110111010110: M1r = 2'b00;
			14'b10110111010110: M1r = 2'b00;
			14'b11110111010110: M1r = 2'b00;
			14'b00001011010110: M1r = 2'b01;
			14'b01001011010110: M1r = 2'b10;
			14'b10001011010110: M1r = 2'b10;
			14'b11001011010110: M1r = 2'b10;
			14'b00011011010110: M1r = 2'b01;
			14'b01011011010110: M1r = 2'b01;
			14'b10011011010110: M1r = 2'b01;
			14'b11011011010110: M1r = 2'b01;
			14'b00101011010110: M1r = 2'b00;
			14'b01101011010110: M1r = 2'b01;
			14'b10101011010110: M1r = 2'b01;
			14'b11101011010110: M1r = 2'b01;
			14'b00111011010110: M1r = 2'b00;
			14'b01111011010110: M1r = 2'b00;
			14'b10111011010110: M1r = 2'b00;
			14'b11111011010110: M1r = 2'b00;
			14'b00001111010110: M1r = 2'b10;
			14'b01001111010110: M1r = 2'b10;
			14'b10001111010110: M1r = 2'b10;
			14'b11001111010110: M1r = 2'b11;
			14'b00011111010110: M1r = 2'b10;
			14'b01011111010110: M1r = 2'b10;
			14'b10011111010110: M1r = 2'b10;
			14'b11011111010110: M1r = 2'b10;
			14'b00101111010110: M1r = 2'b01;
			14'b01101111010110: M1r = 2'b01;
			14'b10101111010110: M1r = 2'b10;
			14'b11101111010110: M1r = 2'b10;
			14'b00111111010110: M1r = 2'b01;
			14'b01111111010110: M1r = 2'b01;
			14'b10111111010110: M1r = 2'b01;
			14'b11111111010110: M1r = 2'b01;
			14'b00000000100110: M1r = 2'b01;
			14'b01000000100110: M1r = 2'b01;
			14'b10000000100110: M1r = 2'b01;
			14'b11000000100110: M1r = 2'b10;
			14'b00010000100110: M1r = 2'b01;
			14'b01010000100110: M1r = 2'b01;
			14'b10010000100110: M1r = 2'b01;
			14'b11010000100110: M1r = 2'b01;
			14'b00100000100110: M1r = 2'b00;
			14'b01100000100110: M1r = 2'b00;
			14'b10100000100110: M1r = 2'b01;
			14'b11100000100110: M1r = 2'b01;
			14'b00110000100110: M1r = 2'b00;
			14'b01110000100110: M1r = 2'b00;
			14'b10110000100110: M1r = 2'b00;
			14'b11110000100110: M1r = 2'b00;
			14'b00000100100110: M1r = 2'b10;
			14'b01000100100110: M1r = 2'b10;
			14'b10000100100110: M1r = 2'b10;
			14'b11000100100110: M1r = 2'b10;
			14'b00010100100110: M1r = 2'b01;
			14'b01010100100110: M1r = 2'b10;
			14'b10010100100110: M1r = 2'b10;
			14'b11010100100110: M1r = 2'b10;
			14'b00100100100110: M1r = 2'b01;
			14'b01100100100110: M1r = 2'b01;
			14'b10100100100110: M1r = 2'b01;
			14'b11100100100110: M1r = 2'b01;
			14'b00110100100110: M1r = 2'b00;
			14'b01110100100110: M1r = 2'b01;
			14'b10110100100110: M1r = 2'b01;
			14'b11110100100110: M1r = 2'b01;
			14'b00001000100110: M1r = 2'b11;
			14'b01001000100110: M1r = 2'b11;
			14'b10001000100110: M1r = 2'b11;
			14'b11001000100110: M1r = 2'b11;
			14'b00011000100110: M1r = 2'b10;
			14'b01011000100110: M1r = 2'b10;
			14'b10011000100110: M1r = 2'b10;
			14'b11011000100110: M1r = 2'b11;
			14'b00101000100110: M1r = 2'b10;
			14'b01101000100110: M1r = 2'b10;
			14'b10101000100110: M1r = 2'b10;
			14'b11101000100110: M1r = 2'b10;
			14'b00111000100110: M1r = 2'b01;
			14'b01111000100110: M1r = 2'b01;
			14'b10111000100110: M1r = 2'b10;
			14'b11111000100110: M1r = 2'b10;
			14'b00001100100110: M1r = 2'b11;
			14'b01001100100110: M1r = 2'b11;
			14'b10001100100110: M1r = 2'b11;
			14'b11001100100110: M1r = 2'b11;
			14'b00011100100110: M1r = 2'b11;
			14'b01011100100110: M1r = 2'b11;
			14'b10011100100110: M1r = 2'b11;
			14'b11011100100110: M1r = 2'b11;
			14'b00101100100110: M1r = 2'b10;
			14'b01101100100110: M1r = 2'b11;
			14'b10101100100110: M1r = 2'b11;
			14'b11101100100110: M1r = 2'b11;
			14'b00111100100110: M1r = 2'b10;
			14'b01111100100110: M1r = 2'b10;
			14'b10111100100110: M1r = 2'b10;
			14'b11111100100110: M1r = 2'b10;
			14'b00000001100110: M1r = 2'b01;
			14'b01000001100110: M1r = 2'b01;
			14'b10000001100110: M1r = 2'b01;
			14'b11000001100110: M1r = 2'b01;
			14'b00010001100110: M1r = 2'b00;
			14'b01010001100110: M1r = 2'b01;
			14'b10010001100110: M1r = 2'b01;
			14'b11010001100110: M1r = 2'b01;
			14'b00100001100110: M1r = 2'b00;
			14'b01100001100110: M1r = 2'b00;
			14'b10100001100110: M1r = 2'b00;
			14'b11100001100110: M1r = 2'b00;
			14'b00110001100110: M1r = 2'b00;
			14'b01110001100110: M1r = 2'b00;
			14'b10110001100110: M1r = 2'b00;
			14'b11110001100110: M1r = 2'b00;
			14'b00000101100110: M1r = 2'b10;
			14'b01000101100110: M1r = 2'b10;
			14'b10000101100110: M1r = 2'b10;
			14'b11000101100110: M1r = 2'b10;
			14'b00010101100110: M1r = 2'b01;
			14'b01010101100110: M1r = 2'b01;
			14'b10010101100110: M1r = 2'b01;
			14'b11010101100110: M1r = 2'b10;
			14'b00100101100110: M1r = 2'b01;
			14'b01100101100110: M1r = 2'b01;
			14'b10100101100110: M1r = 2'b01;
			14'b11100101100110: M1r = 2'b01;
			14'b00110101100110: M1r = 2'b00;
			14'b01110101100110: M1r = 2'b00;
			14'b10110101100110: M1r = 2'b01;
			14'b11110101100110: M1r = 2'b01;
			14'b00001001100110: M1r = 2'b10;
			14'b01001001100110: M1r = 2'b11;
			14'b10001001100110: M1r = 2'b11;
			14'b11001001100110: M1r = 2'b11;
			14'b00011001100110: M1r = 2'b10;
			14'b01011001100110: M1r = 2'b10;
			14'b10011001100110: M1r = 2'b10;
			14'b11011001100110: M1r = 2'b10;
			14'b00101001100110: M1r = 2'b01;
			14'b01101001100110: M1r = 2'b10;
			14'b10101001100110: M1r = 2'b10;
			14'b11101001100110: M1r = 2'b10;
			14'b00111001100110: M1r = 2'b01;
			14'b01111001100110: M1r = 2'b01;
			14'b10111001100110: M1r = 2'b01;
			14'b11111001100110: M1r = 2'b01;
			14'b00001101100110: M1r = 2'b11;
			14'b01001101100110: M1r = 2'b11;
			14'b10001101100110: M1r = 2'b11;
			14'b11001101100110: M1r = 2'b11;
			14'b00011101100110: M1r = 2'b11;
			14'b01011101100110: M1r = 2'b11;
			14'b10011101100110: M1r = 2'b11;
			14'b11011101100110: M1r = 2'b11;
			14'b00101101100110: M1r = 2'b10;
			14'b01101101100110: M1r = 2'b10;
			14'b10101101100110: M1r = 2'b10;
			14'b11101101100110: M1r = 2'b11;
			14'b00111101100110: M1r = 2'b10;
			14'b01111101100110: M1r = 2'b10;
			14'b10111101100110: M1r = 2'b10;
			14'b11111101100110: M1r = 2'b10;
			14'b00000010100110: M1r = 2'b01;
			14'b01000010100110: M1r = 2'b01;
			14'b10000010100110: M1r = 2'b01;
			14'b11000010100110: M1r = 2'b01;
			14'b00010010100110: M1r = 2'b00;
			14'b01010010100110: M1r = 2'b00;
			14'b10010010100110: M1r = 2'b00;
			14'b11010010100110: M1r = 2'b01;
			14'b00100010100110: M1r = 2'b00;
			14'b01100010100110: M1r = 2'b00;
			14'b10100010100110: M1r = 2'b00;
			14'b11100010100110: M1r = 2'b00;
			14'b00110010100110: M1r = 2'b00;
			14'b01110010100110: M1r = 2'b00;
			14'b10110010100110: M1r = 2'b00;
			14'b11110010100110: M1r = 2'b00;
			14'b00000110100110: M1r = 2'b01;
			14'b01000110100110: M1r = 2'b10;
			14'b10000110100110: M1r = 2'b10;
			14'b11000110100110: M1r = 2'b10;
			14'b00010110100110: M1r = 2'b01;
			14'b01010110100110: M1r = 2'b01;
			14'b10010110100110: M1r = 2'b01;
			14'b11010110100110: M1r = 2'b01;
			14'b00100110100110: M1r = 2'b00;
			14'b01100110100110: M1r = 2'b01;
			14'b10100110100110: M1r = 2'b01;
			14'b11100110100110: M1r = 2'b01;
			14'b00110110100110: M1r = 2'b00;
			14'b01110110100110: M1r = 2'b00;
			14'b10110110100110: M1r = 2'b00;
			14'b11110110100110: M1r = 2'b00;
			14'b00001010100110: M1r = 2'b10;
			14'b01001010100110: M1r = 2'b10;
			14'b10001010100110: M1r = 2'b10;
			14'b11001010100110: M1r = 2'b11;
			14'b00011010100110: M1r = 2'b10;
			14'b01011010100110: M1r = 2'b10;
			14'b10011010100110: M1r = 2'b10;
			14'b11011010100110: M1r = 2'b10;
			14'b00101010100110: M1r = 2'b01;
			14'b01101010100110: M1r = 2'b01;
			14'b10101010100110: M1r = 2'b01;
			14'b11101010100110: M1r = 2'b10;
			14'b00111010100110: M1r = 2'b01;
			14'b01111010100110: M1r = 2'b01;
			14'b10111010100110: M1r = 2'b01;
			14'b11111010100110: M1r = 2'b01;
			14'b00001110100110: M1r = 2'b11;
			14'b01001110100110: M1r = 2'b11;
			14'b10001110100110: M1r = 2'b11;
			14'b11001110100110: M1r = 2'b11;
			14'b00011110100110: M1r = 2'b10;
			14'b01011110100110: M1r = 2'b11;
			14'b10011110100110: M1r = 2'b11;
			14'b11011110100110: M1r = 2'b11;
			14'b00101110100110: M1r = 2'b10;
			14'b01101110100110: M1r = 2'b10;
			14'b10101110100110: M1r = 2'b10;
			14'b11101110100110: M1r = 2'b10;
			14'b00111110100110: M1r = 2'b01;
			14'b01111110100110: M1r = 2'b10;
			14'b10111110100110: M1r = 2'b10;
			14'b11111110100110: M1r = 2'b10;
			14'b00000011100110: M1r = 2'b00;
			14'b01000011100110: M1r = 2'b00;
			14'b10000011100110: M1r = 2'b01;
			14'b11000011100110: M1r = 2'b01;
			14'b00010011100110: M1r = 2'b00;
			14'b01010011100110: M1r = 2'b00;
			14'b10010011100110: M1r = 2'b00;
			14'b11010011100110: M1r = 2'b00;
			14'b00100011100110: M1r = 2'b00;
			14'b01100011100110: M1r = 2'b00;
			14'b10100011100110: M1r = 2'b00;
			14'b11100011100110: M1r = 2'b00;
			14'b00110011100110: M1r = 2'b00;
			14'b01110011100110: M1r = 2'b00;
			14'b10110011100110: M1r = 2'b00;
			14'b11110011100110: M1r = 2'b00;
			14'b00000111100110: M1r = 2'b01;
			14'b01000111100110: M1r = 2'b01;
			14'b10000111100110: M1r = 2'b01;
			14'b11000111100110: M1r = 2'b10;
			14'b00010111100110: M1r = 2'b01;
			14'b01010111100110: M1r = 2'b01;
			14'b10010111100110: M1r = 2'b01;
			14'b11010111100110: M1r = 2'b01;
			14'b00100111100110: M1r = 2'b00;
			14'b01100111100110: M1r = 2'b00;
			14'b10100111100110: M1r = 2'b00;
			14'b11100111100110: M1r = 2'b01;
			14'b00110111100110: M1r = 2'b00;
			14'b01110111100110: M1r = 2'b00;
			14'b10110111100110: M1r = 2'b00;
			14'b11110111100110: M1r = 2'b00;
			14'b00001011100110: M1r = 2'b10;
			14'b01001011100110: M1r = 2'b10;
			14'b10001011100110: M1r = 2'b10;
			14'b11001011100110: M1r = 2'b10;
			14'b00011011100110: M1r = 2'b01;
			14'b01011011100110: M1r = 2'b10;
			14'b10011011100110: M1r = 2'b10;
			14'b11011011100110: M1r = 2'b10;
			14'b00101011100110: M1r = 2'b01;
			14'b01101011100110: M1r = 2'b01;
			14'b10101011100110: M1r = 2'b01;
			14'b11101011100110: M1r = 2'b01;
			14'b00111011100110: M1r = 2'b00;
			14'b01111011100110: M1r = 2'b01;
			14'b10111011100110: M1r = 2'b01;
			14'b11111011100110: M1r = 2'b01;
			14'b00001111100110: M1r = 2'b11;
			14'b01001111100110: M1r = 2'b11;
			14'b10001111100110: M1r = 2'b11;
			14'b11001111100110: M1r = 2'b11;
			14'b00011111100110: M1r = 2'b10;
			14'b01011111100110: M1r = 2'b10;
			14'b10011111100110: M1r = 2'b10;
			14'b11011111100110: M1r = 2'b11;
			14'b00101111100110: M1r = 2'b10;
			14'b01101111100110: M1r = 2'b10;
			14'b10101111100110: M1r = 2'b10;
			14'b11101111100110: M1r = 2'b10;
			14'b00111111100110: M1r = 2'b01;
			14'b01111111100110: M1r = 2'b01;
			14'b10111111100110: M1r = 2'b01;
			14'b11111111100110: M1r = 2'b10;
			14'b00000000110110: M1r = 2'b10;
			14'b01000000110110: M1r = 2'b10;
			14'b10000000110110: M1r = 2'b10;
			14'b11000000110110: M1r = 2'b10;
			14'b00010000110110: M1r = 2'b01;
			14'b01010000110110: M1r = 2'b01;
			14'b10010000110110: M1r = 2'b01;
			14'b11010000110110: M1r = 2'b10;
			14'b00100000110110: M1r = 2'b01;
			14'b01100000110110: M1r = 2'b01;
			14'b10100000110110: M1r = 2'b01;
			14'b11100000110110: M1r = 2'b01;
			14'b00110000110110: M1r = 2'b00;
			14'b01110000110110: M1r = 2'b00;
			14'b10110000110110: M1r = 2'b00;
			14'b11110000110110: M1r = 2'b01;
			14'b00000100110110: M1r = 2'b10;
			14'b01000100110110: M1r = 2'b10;
			14'b10000100110110: M1r = 2'b11;
			14'b11000100110110: M1r = 2'b11;
			14'b00010100110110: M1r = 2'b10;
			14'b01010100110110: M1r = 2'b10;
			14'b10010100110110: M1r = 2'b10;
			14'b11010100110110: M1r = 2'b10;
			14'b00100100110110: M1r = 2'b01;
			14'b01100100110110: M1r = 2'b10;
			14'b10100100110110: M1r = 2'b10;
			14'b11100100110110: M1r = 2'b10;
			14'b00110100110110: M1r = 2'b01;
			14'b01110100110110: M1r = 2'b01;
			14'b10110100110110: M1r = 2'b01;
			14'b11110100110110: M1r = 2'b01;
			14'b00001000110110: M1r = 2'b11;
			14'b01001000110110: M1r = 2'b11;
			14'b10001000110110: M1r = 2'b11;
			14'b11001000110110: M1r = 2'b11;
			14'b00011000110110: M1r = 2'b11;
			14'b01011000110110: M1r = 2'b11;
			14'b10011000110110: M1r = 2'b11;
			14'b11011000110110: M1r = 2'b11;
			14'b00101000110110: M1r = 2'b10;
			14'b01101000110110: M1r = 2'b10;
			14'b10101000110110: M1r = 2'b10;
			14'b11101000110110: M1r = 2'b11;
			14'b00111000110110: M1r = 2'b10;
			14'b01111000110110: M1r = 2'b10;
			14'b10111000110110: M1r = 2'b10;
			14'b11111000110110: M1r = 2'b10;
			14'b00001100110110: M1r = 2'b11;
			14'b01001100110110: M1r = 2'b11;
			14'b10001100110110: M1r = 2'b11;
			14'b11001100110110: M1r = 2'b11;
			14'b00011100110110: M1r = 2'b11;
			14'b01011100110110: M1r = 2'b11;
			14'b10011100110110: M1r = 2'b11;
			14'b11011100110110: M1r = 2'b11;
			14'b00101100110110: M1r = 2'b11;
			14'b01101100110110: M1r = 2'b11;
			14'b10101100110110: M1r = 2'b11;
			14'b11101100110110: M1r = 2'b11;
			14'b00111100110110: M1r = 2'b10;
			14'b01111100110110: M1r = 2'b11;
			14'b10111100110110: M1r = 2'b11;
			14'b11111100110110: M1r = 2'b11;
			14'b00000001110110: M1r = 2'b01;
			14'b01000001110110: M1r = 2'b01;
			14'b10000001110110: M1r = 2'b10;
			14'b11000001110110: M1r = 2'b10;
			14'b00010001110110: M1r = 2'b01;
			14'b01010001110110: M1r = 2'b01;
			14'b10010001110110: M1r = 2'b01;
			14'b11010001110110: M1r = 2'b01;
			14'b00100001110110: M1r = 2'b00;
			14'b01100001110110: M1r = 2'b01;
			14'b10100001110110: M1r = 2'b01;
			14'b11100001110110: M1r = 2'b01;
			14'b00110001110110: M1r = 2'b00;
			14'b01110001110110: M1r = 2'b00;
			14'b10110001110110: M1r = 2'b00;
			14'b11110001110110: M1r = 2'b00;
			14'b00000101110110: M1r = 2'b10;
			14'b01000101110110: M1r = 2'b10;
			14'b10000101110110: M1r = 2'b10;
			14'b11000101110110: M1r = 2'b11;
			14'b00010101110110: M1r = 2'b10;
			14'b01010101110110: M1r = 2'b10;
			14'b10010101110110: M1r = 2'b10;
			14'b11010101110110: M1r = 2'b10;
			14'b00100101110110: M1r = 2'b01;
			14'b01100101110110: M1r = 2'b01;
			14'b10100101110110: M1r = 2'b01;
			14'b11100101110110: M1r = 2'b10;
			14'b00110101110110: M1r = 2'b01;
			14'b01110101110110: M1r = 2'b01;
			14'b10110101110110: M1r = 2'b01;
			14'b11110101110110: M1r = 2'b01;
			14'b00001001110110: M1r = 2'b11;
			14'b01001001110110: M1r = 2'b11;
			14'b10001001110110: M1r = 2'b11;
			14'b11001001110110: M1r = 2'b11;
			14'b00011001110110: M1r = 2'b10;
			14'b01011001110110: M1r = 2'b10;
			14'b10011001110110: M1r = 2'b11;
			14'b11011001110110: M1r = 2'b11;
			14'b00101001110110: M1r = 2'b10;
			14'b01101001110110: M1r = 2'b10;
			14'b10101001110110: M1r = 2'b10;
			14'b11101001110110: M1r = 2'b10;
			14'b00111001110110: M1r = 2'b01;
			14'b01111001110110: M1r = 2'b10;
			14'b10111001110110: M1r = 2'b10;
			14'b11111001110110: M1r = 2'b10;
			14'b00001101110110: M1r = 2'b11;
			14'b01001101110110: M1r = 2'b11;
			14'b10001101110110: M1r = 2'b11;
			14'b11001101110110: M1r = 2'b11;
			14'b00011101110110: M1r = 2'b11;
			14'b01011101110110: M1r = 2'b11;
			14'b10011101110110: M1r = 2'b11;
			14'b11011101110110: M1r = 2'b11;
			14'b00101101110110: M1r = 2'b11;
			14'b01101101110110: M1r = 2'b11;
			14'b10101101110110: M1r = 2'b11;
			14'b11101101110110: M1r = 2'b11;
			14'b00111101110110: M1r = 2'b10;
			14'b01111101110110: M1r = 2'b10;
			14'b10111101110110: M1r = 2'b10;
			14'b11111101110110: M1r = 2'b11;
			14'b00000010110110: M1r = 2'b01;
			14'b01000010110110: M1r = 2'b01;
			14'b10000010110110: M1r = 2'b01;
			14'b11000010110110: M1r = 2'b10;
			14'b00010010110110: M1r = 2'b01;
			14'b01010010110110: M1r = 2'b01;
			14'b10010010110110: M1r = 2'b01;
			14'b11010010110110: M1r = 2'b01;
			14'b00100010110110: M1r = 2'b00;
			14'b01100010110110: M1r = 2'b00;
			14'b10100010110110: M1r = 2'b00;
			14'b11100010110110: M1r = 2'b01;
			14'b00110010110110: M1r = 2'b00;
			14'b01110010110110: M1r = 2'b00;
			14'b10110010110110: M1r = 2'b00;
			14'b11110010110110: M1r = 2'b00;
			14'b00000110110110: M1r = 2'b10;
			14'b01000110110110: M1r = 2'b10;
			14'b10000110110110: M1r = 2'b10;
			14'b11000110110110: M1r = 2'b10;
			14'b00010110110110: M1r = 2'b01;
			14'b01010110110110: M1r = 2'b01;
			14'b10010110110110: M1r = 2'b10;
			14'b11010110110110: M1r = 2'b10;
			14'b00100110110110: M1r = 2'b01;
			14'b01100110110110: M1r = 2'b01;
			14'b10100110110110: M1r = 2'b01;
			14'b11100110110110: M1r = 2'b01;
			14'b00110110110110: M1r = 2'b00;
			14'b01110110110110: M1r = 2'b01;
			14'b10110110110110: M1r = 2'b01;
			14'b11110110110110: M1r = 2'b01;
			14'b00001010110110: M1r = 2'b11;
			14'b01001010110110: M1r = 2'b11;
			14'b10001010110110: M1r = 2'b11;
			14'b11001010110110: M1r = 2'b11;
			14'b00011010110110: M1r = 2'b10;
			14'b01011010110110: M1r = 2'b10;
			14'b10011010110110: M1r = 2'b10;
			14'b11011010110110: M1r = 2'b11;
			14'b00101010110110: M1r = 2'b10;
			14'b01101010110110: M1r = 2'b10;
			14'b10101010110110: M1r = 2'b10;
			14'b11101010110110: M1r = 2'b10;
			14'b00111010110110: M1r = 2'b01;
			14'b01111010110110: M1r = 2'b01;
			14'b10111010110110: M1r = 2'b01;
			14'b11111010110110: M1r = 2'b10;
			14'b00001110110110: M1r = 2'b11;
			14'b01001110110110: M1r = 2'b11;
			14'b10001110110110: M1r = 2'b11;
			14'b11001110110110: M1r = 2'b11;
			14'b00011110110110: M1r = 2'b11;
			14'b01011110110110: M1r = 2'b11;
			14'b10011110110110: M1r = 2'b11;
			14'b11011110110110: M1r = 2'b11;
			14'b00101110110110: M1r = 2'b10;
			14'b01101110110110: M1r = 2'b10;
			14'b10101110110110: M1r = 2'b11;
			14'b11101110110110: M1r = 2'b11;
			14'b00111110110110: M1r = 2'b10;
			14'b01111110110110: M1r = 2'b10;
			14'b10111110110110: M1r = 2'b10;
			14'b11111110110110: M1r = 2'b10;
			14'b00000011110110: M1r = 2'b01;
			14'b01000011110110: M1r = 2'b01;
			14'b10000011110110: M1r = 2'b01;
			14'b11000011110110: M1r = 2'b01;
			14'b00010011110110: M1r = 2'b00;
			14'b01010011110110: M1r = 2'b00;
			14'b10010011110110: M1r = 2'b01;
			14'b11010011110110: M1r = 2'b01;
			14'b00100011110110: M1r = 2'b00;
			14'b01100011110110: M1r = 2'b00;
			14'b10100011110110: M1r = 2'b00;
			14'b11100011110110: M1r = 2'b00;
			14'b00110011110110: M1r = 2'b00;
			14'b01110011110110: M1r = 2'b00;
			14'b10110011110110: M1r = 2'b00;
			14'b11110011110110: M1r = 2'b00;
			14'b00000111110110: M1r = 2'b10;
			14'b01000111110110: M1r = 2'b10;
			14'b10000111110110: M1r = 2'b10;
			14'b11000111110110: M1r = 2'b10;
			14'b00010111110110: M1r = 2'b01;
			14'b01010111110110: M1r = 2'b01;
			14'b10010111110110: M1r = 2'b01;
			14'b11010111110110: M1r = 2'b10;
			14'b00100111110110: M1r = 2'b01;
			14'b01100111110110: M1r = 2'b01;
			14'b10100111110110: M1r = 2'b01;
			14'b11100111110110: M1r = 2'b01;
			14'b00110111110110: M1r = 2'b00;
			14'b01110111110110: M1r = 2'b00;
			14'b10110111110110: M1r = 2'b00;
			14'b11110111110110: M1r = 2'b01;
			14'b00001011110110: M1r = 2'b10;
			14'b01001011110110: M1r = 2'b10;
			14'b10001011110110: M1r = 2'b11;
			14'b11001011110110: M1r = 2'b11;
			14'b00011011110110: M1r = 2'b10;
			14'b01011011110110: M1r = 2'b10;
			14'b10011011110110: M1r = 2'b10;
			14'b11011011110110: M1r = 2'b10;
			14'b00101011110110: M1r = 2'b01;
			14'b01101011110110: M1r = 2'b01;
			14'b10101011110110: M1r = 2'b10;
			14'b11101011110110: M1r = 2'b10;
			14'b00111011110110: M1r = 2'b01;
			14'b01111011110110: M1r = 2'b01;
			14'b10111011110110: M1r = 2'b01;
			14'b11111011110110: M1r = 2'b01;
			14'b00001111110110: M1r = 2'b11;
			14'b01001111110110: M1r = 2'b11;
			14'b10001111110110: M1r = 2'b11;
			14'b11001111110110: M1r = 2'b11;
			14'b00011111110110: M1r = 2'b11;
			14'b01011111110110: M1r = 2'b11;
			14'b10011111110110: M1r = 2'b11;
			14'b11011111110110: M1r = 2'b11;
			14'b00101111110110: M1r = 2'b10;
			14'b01101111110110: M1r = 2'b10;
			14'b10101111110110: M1r = 2'b10;
			14'b11101111110110: M1r = 2'b11;
			14'b00111111110110: M1r = 2'b10;
			14'b01111111110110: M1r = 2'b10;
			14'b10111111110110: M1r = 2'b10;
			14'b11111111110110: M1r = 2'b10;
			14'b00000000001010: M1r = 2'b00;
			14'b01000000001010: M1r = 2'b00;
			14'b10000000001010: M1r = 2'b00;
			14'b11000000001010: M1r = 2'b00;
			14'b00010000001010: M1r = 2'b00;
			14'b01010000001010: M1r = 2'b00;
			14'b10010000001010: M1r = 2'b00;
			14'b11010000001010: M1r = 2'b00;
			14'b00100000001010: M1r = 2'b00;
			14'b01100000001010: M1r = 2'b00;
			14'b10100000001010: M1r = 2'b00;
			14'b11100000001010: M1r = 2'b00;
			14'b00110000001010: M1r = 2'b00;
			14'b01110000001010: M1r = 2'b00;
			14'b10110000001010: M1r = 2'b00;
			14'b11110000001010: M1r = 2'b00;
			14'b00000100001010: M1r = 2'b00;
			14'b01000100001010: M1r = 2'b00;
			14'b10000100001010: M1r = 2'b01;
			14'b11000100001010: M1r = 2'b01;
			14'b00010100001010: M1r = 2'b00;
			14'b01010100001010: M1r = 2'b00;
			14'b10010100001010: M1r = 2'b00;
			14'b11010100001010: M1r = 2'b00;
			14'b00100100001010: M1r = 2'b00;
			14'b01100100001010: M1r = 2'b00;
			14'b10100100001010: M1r = 2'b00;
			14'b11100100001010: M1r = 2'b00;
			14'b00110100001010: M1r = 2'b00;
			14'b01110100001010: M1r = 2'b00;
			14'b10110100001010: M1r = 2'b00;
			14'b11110100001010: M1r = 2'b00;
			14'b00001000001010: M1r = 2'b01;
			14'b01001000001010: M1r = 2'b01;
			14'b10001000001010: M1r = 2'b01;
			14'b11001000001010: M1r = 2'b01;
			14'b00011000001010: M1r = 2'b01;
			14'b01011000001010: M1r = 2'b01;
			14'b10011000001010: M1r = 2'b01;
			14'b11011000001010: M1r = 2'b01;
			14'b00101000001010: M1r = 2'b00;
			14'b01101000001010: M1r = 2'b00;
			14'b10101000001010: M1r = 2'b00;
			14'b11101000001010: M1r = 2'b01;
			14'b00111000001010: M1r = 2'b00;
			14'b01111000001010: M1r = 2'b00;
			14'b10111000001010: M1r = 2'b00;
			14'b11111000001010: M1r = 2'b00;
			14'b00001100001010: M1r = 2'b10;
			14'b01001100001010: M1r = 2'b10;
			14'b10001100001010: M1r = 2'b10;
			14'b11001100001010: M1r = 2'b10;
			14'b00011100001010: M1r = 2'b01;
			14'b01011100001010: M1r = 2'b01;
			14'b10011100001010: M1r = 2'b10;
			14'b11011100001010: M1r = 2'b10;
			14'b00101100001010: M1r = 2'b01;
			14'b01101100001010: M1r = 2'b01;
			14'b10101100001010: M1r = 2'b01;
			14'b11101100001010: M1r = 2'b01;
			14'b00111100001010: M1r = 2'b00;
			14'b01111100001010: M1r = 2'b01;
			14'b10111100001010: M1r = 2'b01;
			14'b11111100001010: M1r = 2'b01;
			14'b00000001001010: M1r = 2'b00;
			14'b01000001001010: M1r = 2'b00;
			14'b10000001001010: M1r = 2'b00;
			14'b11000001001010: M1r = 2'b00;
			14'b00010001001010: M1r = 2'b00;
			14'b01010001001010: M1r = 2'b00;
			14'b10010001001010: M1r = 2'b00;
			14'b11010001001010: M1r = 2'b00;
			14'b00100001001010: M1r = 2'b00;
			14'b01100001001010: M1r = 2'b00;
			14'b10100001001010: M1r = 2'b00;
			14'b11100001001010: M1r = 2'b00;
			14'b00110001001010: M1r = 2'b00;
			14'b01110001001010: M1r = 2'b00;
			14'b10110001001010: M1r = 2'b00;
			14'b11110001001010: M1r = 2'b00;
			14'b00000101001010: M1r = 2'b00;
			14'b01000101001010: M1r = 2'b00;
			14'b10000101001010: M1r = 2'b00;
			14'b11000101001010: M1r = 2'b00;
			14'b00010101001010: M1r = 2'b00;
			14'b01010101001010: M1r = 2'b00;
			14'b10010101001010: M1r = 2'b00;
			14'b11010101001010: M1r = 2'b00;
			14'b00100101001010: M1r = 2'b00;
			14'b01100101001010: M1r = 2'b00;
			14'b10100101001010: M1r = 2'b00;
			14'b11100101001010: M1r = 2'b00;
			14'b00110101001010: M1r = 2'b00;
			14'b01110101001010: M1r = 2'b00;
			14'b10110101001010: M1r = 2'b00;
			14'b11110101001010: M1r = 2'b00;
			14'b00001001001010: M1r = 2'b01;
			14'b01001001001010: M1r = 2'b01;
			14'b10001001001010: M1r = 2'b01;
			14'b11001001001010: M1r = 2'b01;
			14'b00011001001010: M1r = 2'b00;
			14'b01011001001010: M1r = 2'b00;
			14'b10011001001010: M1r = 2'b01;
			14'b11011001001010: M1r = 2'b01;
			14'b00101001001010: M1r = 2'b00;
			14'b01101001001010: M1r = 2'b00;
			14'b10101001001010: M1r = 2'b00;
			14'b11101001001010: M1r = 2'b00;
			14'b00111001001010: M1r = 2'b00;
			14'b01111001001010: M1r = 2'b00;
			14'b10111001001010: M1r = 2'b00;
			14'b11111001001010: M1r = 2'b00;
			14'b00001101001010: M1r = 2'b01;
			14'b01001101001010: M1r = 2'b10;
			14'b10001101001010: M1r = 2'b10;
			14'b11001101001010: M1r = 2'b10;
			14'b00011101001010: M1r = 2'b01;
			14'b01011101001010: M1r = 2'b01;
			14'b10011101001010: M1r = 2'b01;
			14'b11011101001010: M1r = 2'b01;
			14'b00101101001010: M1r = 2'b01;
			14'b01101101001010: M1r = 2'b01;
			14'b10101101001010: M1r = 2'b01;
			14'b11101101001010: M1r = 2'b01;
			14'b00111101001010: M1r = 2'b00;
			14'b01111101001010: M1r = 2'b00;
			14'b10111101001010: M1r = 2'b00;
			14'b11111101001010: M1r = 2'b01;
			14'b00000010001010: M1r = 2'b00;
			14'b01000010001010: M1r = 2'b00;
			14'b10000010001010: M1r = 2'b00;
			14'b11000010001010: M1r = 2'b00;
			14'b00010010001010: M1r = 2'b00;
			14'b01010010001010: M1r = 2'b00;
			14'b10010010001010: M1r = 2'b00;
			14'b11010010001010: M1r = 2'b00;
			14'b00100010001010: M1r = 2'b00;
			14'b01100010001010: M1r = 2'b00;
			14'b10100010001010: M1r = 2'b00;
			14'b11100010001010: M1r = 2'b00;
			14'b00110010001010: M1r = 2'b00;
			14'b01110010001010: M1r = 2'b00;
			14'b10110010001010: M1r = 2'b00;
			14'b11110010001010: M1r = 2'b00;
			14'b00000110001010: M1r = 2'b00;
			14'b01000110001010: M1r = 2'b00;
			14'b10000110001010: M1r = 2'b00;
			14'b11000110001010: M1r = 2'b00;
			14'b00010110001010: M1r = 2'b00;
			14'b01010110001010: M1r = 2'b00;
			14'b10010110001010: M1r = 2'b00;
			14'b11010110001010: M1r = 2'b00;
			14'b00100110001010: M1r = 2'b00;
			14'b01100110001010: M1r = 2'b00;
			14'b10100110001010: M1r = 2'b00;
			14'b11100110001010: M1r = 2'b00;
			14'b00110110001010: M1r = 2'b00;
			14'b01110110001010: M1r = 2'b00;
			14'b10110110001010: M1r = 2'b00;
			14'b11110110001010: M1r = 2'b00;
			14'b00001010001010: M1r = 2'b00;
			14'b01001010001010: M1r = 2'b01;
			14'b10001010001010: M1r = 2'b01;
			14'b11001010001010: M1r = 2'b01;
			14'b00011010001010: M1r = 2'b00;
			14'b01011010001010: M1r = 2'b00;
			14'b10011010001010: M1r = 2'b00;
			14'b11011010001010: M1r = 2'b00;
			14'b00101010001010: M1r = 2'b00;
			14'b01101010001010: M1r = 2'b00;
			14'b10101010001010: M1r = 2'b00;
			14'b11101010001010: M1r = 2'b00;
			14'b00111010001010: M1r = 2'b00;
			14'b01111010001010: M1r = 2'b00;
			14'b10111010001010: M1r = 2'b00;
			14'b11111010001010: M1r = 2'b00;
			14'b00001110001010: M1r = 2'b01;
			14'b01001110001010: M1r = 2'b01;
			14'b10001110001010: M1r = 2'b10;
			14'b11001110001010: M1r = 2'b10;
			14'b00011110001010: M1r = 2'b01;
			14'b01011110001010: M1r = 2'b01;
			14'b10011110001010: M1r = 2'b01;
			14'b11011110001010: M1r = 2'b01;
			14'b00101110001010: M1r = 2'b00;
			14'b01101110001010: M1r = 2'b00;
			14'b10101110001010: M1r = 2'b01;
			14'b11101110001010: M1r = 2'b01;
			14'b00111110001010: M1r = 2'b00;
			14'b01111110001010: M1r = 2'b00;
			14'b10111110001010: M1r = 2'b00;
			14'b11111110001010: M1r = 2'b00;
			14'b00000011001010: M1r = 2'b00;
			14'b01000011001010: M1r = 2'b00;
			14'b10000011001010: M1r = 2'b00;
			14'b11000011001010: M1r = 2'b00;
			14'b00010011001010: M1r = 2'b00;
			14'b01010011001010: M1r = 2'b00;
			14'b10010011001010: M1r = 2'b00;
			14'b11010011001010: M1r = 2'b00;
			14'b00100011001010: M1r = 2'b00;
			14'b01100011001010: M1r = 2'b00;
			14'b10100011001010: M1r = 2'b00;
			14'b11100011001010: M1r = 2'b00;
			14'b00110011001010: M1r = 2'b00;
			14'b01110011001010: M1r = 2'b00;
			14'b10110011001010: M1r = 2'b00;
			14'b11110011001010: M1r = 2'b00;
			14'b00000111001010: M1r = 2'b00;
			14'b01000111001010: M1r = 2'b00;
			14'b10000111001010: M1r = 2'b00;
			14'b11000111001010: M1r = 2'b00;
			14'b00010111001010: M1r = 2'b00;
			14'b01010111001010: M1r = 2'b00;
			14'b10010111001010: M1r = 2'b00;
			14'b11010111001010: M1r = 2'b00;
			14'b00100111001010: M1r = 2'b00;
			14'b01100111001010: M1r = 2'b00;
			14'b10100111001010: M1r = 2'b00;
			14'b11100111001010: M1r = 2'b00;
			14'b00110111001010: M1r = 2'b00;
			14'b01110111001010: M1r = 2'b00;
			14'b10110111001010: M1r = 2'b00;
			14'b11110111001010: M1r = 2'b00;
			14'b00001011001010: M1r = 2'b00;
			14'b01001011001010: M1r = 2'b00;
			14'b10001011001010: M1r = 2'b01;
			14'b11001011001010: M1r = 2'b01;
			14'b00011011001010: M1r = 2'b00;
			14'b01011011001010: M1r = 2'b00;
			14'b10011011001010: M1r = 2'b00;
			14'b11011011001010: M1r = 2'b00;
			14'b00101011001010: M1r = 2'b00;
			14'b01101011001010: M1r = 2'b00;
			14'b10101011001010: M1r = 2'b00;
			14'b11101011001010: M1r = 2'b00;
			14'b00111011001010: M1r = 2'b00;
			14'b01111011001010: M1r = 2'b00;
			14'b10111011001010: M1r = 2'b00;
			14'b11111011001010: M1r = 2'b00;
			14'b00001111001010: M1r = 2'b01;
			14'b01001111001010: M1r = 2'b01;
			14'b10001111001010: M1r = 2'b01;
			14'b11001111001010: M1r = 2'b01;
			14'b00011111001010: M1r = 2'b00;
			14'b01011111001010: M1r = 2'b01;
			14'b10011111001010: M1r = 2'b01;
			14'b11011111001010: M1r = 2'b01;
			14'b00101111001010: M1r = 2'b00;
			14'b01101111001010: M1r = 2'b00;
			14'b10101111001010: M1r = 2'b00;
			14'b11101111001010: M1r = 2'b00;
			14'b00111111001010: M1r = 2'b00;
			14'b01111111001010: M1r = 2'b00;
			14'b10111111001010: M1r = 2'b00;
			14'b11111111001010: M1r = 2'b00;
			14'b00000000011010: M1r = 2'b00;
			14'b01000000011010: M1r = 2'b00;
			14'b10000000011010: M1r = 2'b00;
			14'b11000000011010: M1r = 2'b00;
			14'b00010000011010: M1r = 2'b00;
			14'b01010000011010: M1r = 2'b00;
			14'b10010000011010: M1r = 2'b00;
			14'b11010000011010: M1r = 2'b00;
			14'b00100000011010: M1r = 2'b00;
			14'b01100000011010: M1r = 2'b00;
			14'b10100000011010: M1r = 2'b00;
			14'b11100000011010: M1r = 2'b00;
			14'b00110000011010: M1r = 2'b00;
			14'b01110000011010: M1r = 2'b00;
			14'b10110000011010: M1r = 2'b00;
			14'b11110000011010: M1r = 2'b00;
			14'b00000100011010: M1r = 2'b01;
			14'b01000100011010: M1r = 2'b01;
			14'b10000100011010: M1r = 2'b01;
			14'b11000100011010: M1r = 2'b01;
			14'b00010100011010: M1r = 2'b00;
			14'b01010100011010: M1r = 2'b00;
			14'b10010100011010: M1r = 2'b01;
			14'b11010100011010: M1r = 2'b01;
			14'b00100100011010: M1r = 2'b00;
			14'b01100100011010: M1r = 2'b00;
			14'b10100100011010: M1r = 2'b00;
			14'b11100100011010: M1r = 2'b00;
			14'b00110100011010: M1r = 2'b00;
			14'b01110100011010: M1r = 2'b00;
			14'b10110100011010: M1r = 2'b00;
			14'b11110100011010: M1r = 2'b00;
			14'b00001000011010: M1r = 2'b01;
			14'b01001000011010: M1r = 2'b10;
			14'b10001000011010: M1r = 2'b10;
			14'b11001000011010: M1r = 2'b10;
			14'b00011000011010: M1r = 2'b01;
			14'b01011000011010: M1r = 2'b01;
			14'b10011000011010: M1r = 2'b01;
			14'b11011000011010: M1r = 2'b01;
			14'b00101000011010: M1r = 2'b01;
			14'b01101000011010: M1r = 2'b01;
			14'b10101000011010: M1r = 2'b01;
			14'b11101000011010: M1r = 2'b01;
			14'b00111000011010: M1r = 2'b00;
			14'b01111000011010: M1r = 2'b00;
			14'b10111000011010: M1r = 2'b00;
			14'b11111000011010: M1r = 2'b00;
			14'b00001100011010: M1r = 2'b10;
			14'b01001100011010: M1r = 2'b10;
			14'b10001100011010: M1r = 2'b11;
			14'b11001100011010: M1r = 2'b11;
			14'b00011100011010: M1r = 2'b10;
			14'b01011100011010: M1r = 2'b10;
			14'b10011100011010: M1r = 2'b10;
			14'b11011100011010: M1r = 2'b10;
			14'b00101100011010: M1r = 2'b01;
			14'b01101100011010: M1r = 2'b01;
			14'b10101100011010: M1r = 2'b10;
			14'b11101100011010: M1r = 2'b10;
			14'b00111100011010: M1r = 2'b01;
			14'b01111100011010: M1r = 2'b01;
			14'b10111100011010: M1r = 2'b01;
			14'b11111100011010: M1r = 2'b01;
			14'b00000001011010: M1r = 2'b00;
			14'b01000001011010: M1r = 2'b00;
			14'b10000001011010: M1r = 2'b00;
			14'b11000001011010: M1r = 2'b00;
			14'b00010001011010: M1r = 2'b00;
			14'b01010001011010: M1r = 2'b00;
			14'b10010001011010: M1r = 2'b00;
			14'b11010001011010: M1r = 2'b00;
			14'b00100001011010: M1r = 2'b00;
			14'b01100001011010: M1r = 2'b00;
			14'b10100001011010: M1r = 2'b00;
			14'b11100001011010: M1r = 2'b00;
			14'b00110001011010: M1r = 2'b00;
			14'b01110001011010: M1r = 2'b00;
			14'b10110001011010: M1r = 2'b00;
			14'b11110001011010: M1r = 2'b00;
			14'b00000101011010: M1r = 2'b00;
			14'b01000101011010: M1r = 2'b01;
			14'b10000101011010: M1r = 2'b01;
			14'b11000101011010: M1r = 2'b01;
			14'b00010101011010: M1r = 2'b00;
			14'b01010101011010: M1r = 2'b00;
			14'b10010101011010: M1r = 2'b00;
			14'b11010101011010: M1r = 2'b00;
			14'b00100101011010: M1r = 2'b00;
			14'b01100101011010: M1r = 2'b00;
			14'b10100101011010: M1r = 2'b00;
			14'b11100101011010: M1r = 2'b00;
			14'b00110101011010: M1r = 2'b00;
			14'b01110101011010: M1r = 2'b00;
			14'b10110101011010: M1r = 2'b00;
			14'b11110101011010: M1r = 2'b00;
			14'b00001001011010: M1r = 2'b01;
			14'b01001001011010: M1r = 2'b01;
			14'b10001001011010: M1r = 2'b01;
			14'b11001001011010: M1r = 2'b10;
			14'b00011001011010: M1r = 2'b01;
			14'b01011001011010: M1r = 2'b01;
			14'b10011001011010: M1r = 2'b01;
			14'b11011001011010: M1r = 2'b01;
			14'b00101001011010: M1r = 2'b00;
			14'b01101001011010: M1r = 2'b00;
			14'b10101001011010: M1r = 2'b01;
			14'b11101001011010: M1r = 2'b01;
			14'b00111001011010: M1r = 2'b00;
			14'b01111001011010: M1r = 2'b00;
			14'b10111001011010: M1r = 2'b00;
			14'b11111001011010: M1r = 2'b00;
			14'b00001101011010: M1r = 2'b10;
			14'b01001101011010: M1r = 2'b10;
			14'b10001101011010: M1r = 2'b10;
			14'b11001101011010: M1r = 2'b10;
			14'b00011101011010: M1r = 2'b01;
			14'b01011101011010: M1r = 2'b10;
			14'b10011101011010: M1r = 2'b10;
			14'b11011101011010: M1r = 2'b10;
			14'b00101101011010: M1r = 2'b01;
			14'b01101101011010: M1r = 2'b01;
			14'b10101101011010: M1r = 2'b01;
			14'b11101101011010: M1r = 2'b01;
			14'b00111101011010: M1r = 2'b01;
			14'b01111101011010: M1r = 2'b01;
			14'b10111101011010: M1r = 2'b01;
			14'b11111101011010: M1r = 2'b01;
			14'b00000010011010: M1r = 2'b00;
			14'b01000010011010: M1r = 2'b00;
			14'b10000010011010: M1r = 2'b00;
			14'b11000010011010: M1r = 2'b00;
			14'b00010010011010: M1r = 2'b00;
			14'b01010010011010: M1r = 2'b00;
			14'b10010010011010: M1r = 2'b00;
			14'b11010010011010: M1r = 2'b00;
			14'b00100010011010: M1r = 2'b00;
			14'b01100010011010: M1r = 2'b00;
			14'b10100010011010: M1r = 2'b00;
			14'b11100010011010: M1r = 2'b00;
			14'b00110010011010: M1r = 2'b00;
			14'b01110010011010: M1r = 2'b00;
			14'b10110010011010: M1r = 2'b00;
			14'b11110010011010: M1r = 2'b00;
			14'b00000110011010: M1r = 2'b00;
			14'b01000110011010: M1r = 2'b00;
			14'b10000110011010: M1r = 2'b00;
			14'b11000110011010: M1r = 2'b01;
			14'b00010110011010: M1r = 2'b00;
			14'b01010110011010: M1r = 2'b00;
			14'b10010110011010: M1r = 2'b00;
			14'b11010110011010: M1r = 2'b00;
			14'b00100110011010: M1r = 2'b00;
			14'b01100110011010: M1r = 2'b00;
			14'b10100110011010: M1r = 2'b00;
			14'b11100110011010: M1r = 2'b00;
			14'b00110110011010: M1r = 2'b00;
			14'b01110110011010: M1r = 2'b00;
			14'b10110110011010: M1r = 2'b00;
			14'b11110110011010: M1r = 2'b00;
			14'b00001010011010: M1r = 2'b01;
			14'b01001010011010: M1r = 2'b01;
			14'b10001010011010: M1r = 2'b01;
			14'b11001010011010: M1r = 2'b01;
			14'b00011010011010: M1r = 2'b00;
			14'b01011010011010: M1r = 2'b01;
			14'b10011010011010: M1r = 2'b01;
			14'b11011010011010: M1r = 2'b01;
			14'b00101010011010: M1r = 2'b00;
			14'b01101010011010: M1r = 2'b00;
			14'b10101010011010: M1r = 2'b00;
			14'b11101010011010: M1r = 2'b00;
			14'b00111010011010: M1r = 2'b00;
			14'b01111010011010: M1r = 2'b00;
			14'b10111010011010: M1r = 2'b00;
			14'b11111010011010: M1r = 2'b00;
			14'b00001110011010: M1r = 2'b10;
			14'b01001110011010: M1r = 2'b10;
			14'b10001110011010: M1r = 2'b10;
			14'b11001110011010: M1r = 2'b10;
			14'b00011110011010: M1r = 2'b01;
			14'b01011110011010: M1r = 2'b01;
			14'b10011110011010: M1r = 2'b01;
			14'b11011110011010: M1r = 2'b10;
			14'b00101110011010: M1r = 2'b01;
			14'b01101110011010: M1r = 2'b01;
			14'b10101110011010: M1r = 2'b01;
			14'b11101110011010: M1r = 2'b01;
			14'b00111110011010: M1r = 2'b00;
			14'b01111110011010: M1r = 2'b00;
			14'b10111110011010: M1r = 2'b01;
			14'b11111110011010: M1r = 2'b01;
			14'b00000011011010: M1r = 2'b00;
			14'b01000011011010: M1r = 2'b00;
			14'b10000011011010: M1r = 2'b00;
			14'b11000011011010: M1r = 2'b00;
			14'b00010011011010: M1r = 2'b00;
			14'b01010011011010: M1r = 2'b00;
			14'b10010011011010: M1r = 2'b00;
			14'b11010011011010: M1r = 2'b00;
			14'b00100011011010: M1r = 2'b00;
			14'b01100011011010: M1r = 2'b00;
			14'b10100011011010: M1r = 2'b00;
			14'b11100011011010: M1r = 2'b00;
			14'b00110011011010: M1r = 2'b00;
			14'b01110011011010: M1r = 2'b00;
			14'b10110011011010: M1r = 2'b00;
			14'b11110011011010: M1r = 2'b00;
			14'b00000111011010: M1r = 2'b00;
			14'b01000111011010: M1r = 2'b00;
			14'b10000111011010: M1r = 2'b00;
			14'b11000111011010: M1r = 2'b00;
			14'b00010111011010: M1r = 2'b00;
			14'b01010111011010: M1r = 2'b00;
			14'b10010111011010: M1r = 2'b00;
			14'b11010111011010: M1r = 2'b00;
			14'b00100111011010: M1r = 2'b00;
			14'b01100111011010: M1r = 2'b00;
			14'b10100111011010: M1r = 2'b00;
			14'b11100111011010: M1r = 2'b00;
			14'b00110111011010: M1r = 2'b00;
			14'b01110111011010: M1r = 2'b00;
			14'b10110111011010: M1r = 2'b00;
			14'b11110111011010: M1r = 2'b00;
			14'b00001011011010: M1r = 2'b01;
			14'b01001011011010: M1r = 2'b01;
			14'b10001011011010: M1r = 2'b01;
			14'b11001011011010: M1r = 2'b01;
			14'b00011011011010: M1r = 2'b00;
			14'b01011011011010: M1r = 2'b00;
			14'b10011011011010: M1r = 2'b00;
			14'b11011011011010: M1r = 2'b01;
			14'b00101011011010: M1r = 2'b00;
			14'b01101011011010: M1r = 2'b00;
			14'b10101011011010: M1r = 2'b00;
			14'b11101011011010: M1r = 2'b00;
			14'b00111011011010: M1r = 2'b00;
			14'b01111011011010: M1r = 2'b00;
			14'b10111011011010: M1r = 2'b00;
			14'b11111011011010: M1r = 2'b00;
			14'b00001111011010: M1r = 2'b01;
			14'b01001111011010: M1r = 2'b10;
			14'b10001111011010: M1r = 2'b10;
			14'b11001111011010: M1r = 2'b10;
			14'b00011111011010: M1r = 2'b01;
			14'b01011111011010: M1r = 2'b01;
			14'b10011111011010: M1r = 2'b01;
			14'b11011111011010: M1r = 2'b01;
			14'b00101111011010: M1r = 2'b00;
			14'b01101111011010: M1r = 2'b01;
			14'b10101111011010: M1r = 2'b01;
			14'b11101111011010: M1r = 2'b01;
			14'b00111111011010: M1r = 2'b00;
			14'b01111111011010: M1r = 2'b00;
			14'b10111111011010: M1r = 2'b00;
			14'b11111111011010: M1r = 2'b00;
			14'b00000000101010: M1r = 2'b00;
			14'b01000000101010: M1r = 2'b01;
			14'b10000000101010: M1r = 2'b01;
			14'b11000000101010: M1r = 2'b01;
			14'b00010000101010: M1r = 2'b00;
			14'b01010000101010: M1r = 2'b00;
			14'b10010000101010: M1r = 2'b00;
			14'b11010000101010: M1r = 2'b00;
			14'b00100000101010: M1r = 2'b00;
			14'b01100000101010: M1r = 2'b00;
			14'b10100000101010: M1r = 2'b00;
			14'b11100000101010: M1r = 2'b00;
			14'b00110000101010: M1r = 2'b00;
			14'b01110000101010: M1r = 2'b00;
			14'b10110000101010: M1r = 2'b00;
			14'b11110000101010: M1r = 2'b00;
			14'b00000100101010: M1r = 2'b01;
			14'b01000100101010: M1r = 2'b01;
			14'b10000100101010: M1r = 2'b01;
			14'b11000100101010: M1r = 2'b10;
			14'b00010100101010: M1r = 2'b01;
			14'b01010100101010: M1r = 2'b01;
			14'b10010100101010: M1r = 2'b01;
			14'b11010100101010: M1r = 2'b01;
			14'b00100100101010: M1r = 2'b00;
			14'b01100100101010: M1r = 2'b00;
			14'b10100100101010: M1r = 2'b00;
			14'b11100100101010: M1r = 2'b01;
			14'b00110100101010: M1r = 2'b00;
			14'b01110100101010: M1r = 2'b00;
			14'b10110100101010: M1r = 2'b00;
			14'b11110100101010: M1r = 2'b00;
			14'b00001000101010: M1r = 2'b10;
			14'b01001000101010: M1r = 2'b10;
			14'b10001000101010: M1r = 2'b10;
			14'b11001000101010: M1r = 2'b10;
			14'b00011000101010: M1r = 2'b01;
			14'b01011000101010: M1r = 2'b10;
			14'b10011000101010: M1r = 2'b10;
			14'b11011000101010: M1r = 2'b10;
			14'b00101000101010: M1r = 2'b01;
			14'b01101000101010: M1r = 2'b01;
			14'b10101000101010: M1r = 2'b01;
			14'b11101000101010: M1r = 2'b01;
			14'b00111000101010: M1r = 2'b00;
			14'b01111000101010: M1r = 2'b01;
			14'b10111000101010: M1r = 2'b01;
			14'b11111000101010: M1r = 2'b01;
			14'b00001100101010: M1r = 2'b11;
			14'b01001100101010: M1r = 2'b11;
			14'b10001100101010: M1r = 2'b11;
			14'b11001100101010: M1r = 2'b11;
			14'b00011100101010: M1r = 2'b10;
			14'b01011100101010: M1r = 2'b10;
			14'b10011100101010: M1r = 2'b10;
			14'b11011100101010: M1r = 2'b11;
			14'b00101100101010: M1r = 2'b10;
			14'b01101100101010: M1r = 2'b10;
			14'b10101100101010: M1r = 2'b10;
			14'b11101100101010: M1r = 2'b10;
			14'b00111100101010: M1r = 2'b01;
			14'b01111100101010: M1r = 2'b01;
			14'b10111100101010: M1r = 2'b10;
			14'b11111100101010: M1r = 2'b10;
			14'b00000001101010: M1r = 2'b00;
			14'b01000001101010: M1r = 2'b00;
			14'b10000001101010: M1r = 2'b00;
			14'b11000001101010: M1r = 2'b01;
			14'b00010001101010: M1r = 2'b00;
			14'b01010001101010: M1r = 2'b00;
			14'b10010001101010: M1r = 2'b00;
			14'b11010001101010: M1r = 2'b00;
			14'b00100001101010: M1r = 2'b00;
			14'b01100001101010: M1r = 2'b00;
			14'b10100001101010: M1r = 2'b00;
			14'b11100001101010: M1r = 2'b00;
			14'b00110001101010: M1r = 2'b00;
			14'b01110001101010: M1r = 2'b00;
			14'b10110001101010: M1r = 2'b00;
			14'b11110001101010: M1r = 2'b00;
			14'b00000101101010: M1r = 2'b01;
			14'b01000101101010: M1r = 2'b01;
			14'b10000101101010: M1r = 2'b01;
			14'b11000101101010: M1r = 2'b01;
			14'b00010101101010: M1r = 2'b00;
			14'b01010101101010: M1r = 2'b01;
			14'b10010101101010: M1r = 2'b01;
			14'b11010101101010: M1r = 2'b01;
			14'b00100101101010: M1r = 2'b00;
			14'b01100101101010: M1r = 2'b00;
			14'b10100101101010: M1r = 2'b00;
			14'b11100101101010: M1r = 2'b00;
			14'b00110101101010: M1r = 2'b00;
			14'b01110101101010: M1r = 2'b00;
			14'b10110101101010: M1r = 2'b00;
			14'b11110101101010: M1r = 2'b00;
			14'b00001001101010: M1r = 2'b10;
			14'b01001001101010: M1r = 2'b10;
			14'b10001001101010: M1r = 2'b10;
			14'b11001001101010: M1r = 2'b10;
			14'b00011001101010: M1r = 2'b01;
			14'b01011001101010: M1r = 2'b01;
			14'b10011001101010: M1r = 2'b01;
			14'b11011001101010: M1r = 2'b10;
			14'b00101001101010: M1r = 2'b01;
			14'b01101001101010: M1r = 2'b01;
			14'b10101001101010: M1r = 2'b01;
			14'b11101001101010: M1r = 2'b01;
			14'b00111001101010: M1r = 2'b00;
			14'b01111001101010: M1r = 2'b00;
			14'b10111001101010: M1r = 2'b00;
			14'b11111001101010: M1r = 2'b01;
			14'b00001101101010: M1r = 2'b10;
			14'b01001101101010: M1r = 2'b11;
			14'b10001101101010: M1r = 2'b11;
			14'b11001101101010: M1r = 2'b11;
			14'b00011101101010: M1r = 2'b10;
			14'b01011101101010: M1r = 2'b10;
			14'b10011101101010: M1r = 2'b10;
			14'b11011101101010: M1r = 2'b10;
			14'b00101101101010: M1r = 2'b01;
			14'b01101101101010: M1r = 2'b10;
			14'b10101101101010: M1r = 2'b10;
			14'b11101101101010: M1r = 2'b10;
			14'b00111101101010: M1r = 2'b01;
			14'b01111101101010: M1r = 2'b01;
			14'b10111101101010: M1r = 2'b01;
			14'b11111101101010: M1r = 2'b01;
			14'b00000010101010: M1r = 2'b00;
			14'b01000010101010: M1r = 2'b00;
			14'b10000010101010: M1r = 2'b00;
			14'b11000010101010: M1r = 2'b00;
			14'b00010010101010: M1r = 2'b00;
			14'b01010010101010: M1r = 2'b00;
			14'b10010010101010: M1r = 2'b00;
			14'b11010010101010: M1r = 2'b00;
			14'b00100010101010: M1r = 2'b00;
			14'b01100010101010: M1r = 2'b00;
			14'b10100010101010: M1r = 2'b00;
			14'b11100010101010: M1r = 2'b00;
			14'b00110010101010: M1r = 2'b00;
			14'b01110010101010: M1r = 2'b00;
			14'b10110010101010: M1r = 2'b00;
			14'b11110010101010: M1r = 2'b00;
			14'b00000110101010: M1r = 2'b01;
			14'b01000110101010: M1r = 2'b01;
			14'b10000110101010: M1r = 2'b01;
			14'b11000110101010: M1r = 2'b01;
			14'b00010110101010: M1r = 2'b00;
			14'b01010110101010: M1r = 2'b00;
			14'b10010110101010: M1r = 2'b00;
			14'b11010110101010: M1r = 2'b01;
			14'b00100110101010: M1r = 2'b00;
			14'b01100110101010: M1r = 2'b00;
			14'b10100110101010: M1r = 2'b00;
			14'b11100110101010: M1r = 2'b00;
			14'b00110110101010: M1r = 2'b00;
			14'b01110110101010: M1r = 2'b00;
			14'b10110110101010: M1r = 2'b00;
			14'b11110110101010: M1r = 2'b00;
			14'b00001010101010: M1r = 2'b01;
			14'b01001010101010: M1r = 2'b01;
			14'b10001010101010: M1r = 2'b10;
			14'b11001010101010: M1r = 2'b10;
			14'b00011010101010: M1r = 2'b01;
			14'b01011010101010: M1r = 2'b01;
			14'b10011010101010: M1r = 2'b01;
			14'b11011010101010: M1r = 2'b01;
			14'b00101010101010: M1r = 2'b00;
			14'b01101010101010: M1r = 2'b01;
			14'b10101010101010: M1r = 2'b01;
			14'b11101010101010: M1r = 2'b01;
			14'b00111010101010: M1r = 2'b00;
			14'b01111010101010: M1r = 2'b00;
			14'b10111010101010: M1r = 2'b00;
			14'b11111010101010: M1r = 2'b00;
			14'b00001110101010: M1r = 2'b10;
			14'b01001110101010: M1r = 2'b10;
			14'b10001110101010: M1r = 2'b10;
			14'b11001110101010: M1r = 2'b11;
			14'b00011110101010: M1r = 2'b10;
			14'b01011110101010: M1r = 2'b10;
			14'b10011110101010: M1r = 2'b10;
			14'b11011110101010: M1r = 2'b10;
			14'b00101110101010: M1r = 2'b01;
			14'b01101110101010: M1r = 2'b01;
			14'b10101110101010: M1r = 2'b01;
			14'b11101110101010: M1r = 2'b10;
			14'b00111110101010: M1r = 2'b01;
			14'b01111110101010: M1r = 2'b01;
			14'b10111110101010: M1r = 2'b01;
			14'b11111110101010: M1r = 2'b01;
			14'b00000011101010: M1r = 2'b00;
			14'b01000011101010: M1r = 2'b00;
			14'b10000011101010: M1r = 2'b00;
			14'b11000011101010: M1r = 2'b00;
			14'b00010011101010: M1r = 2'b00;
			14'b01010011101010: M1r = 2'b00;
			14'b10010011101010: M1r = 2'b00;
			14'b11010011101010: M1r = 2'b00;
			14'b00100011101010: M1r = 2'b00;
			14'b01100011101010: M1r = 2'b00;
			14'b10100011101010: M1r = 2'b00;
			14'b11100011101010: M1r = 2'b00;
			14'b00110011101010: M1r = 2'b00;
			14'b01110011101010: M1r = 2'b00;
			14'b10110011101010: M1r = 2'b00;
			14'b11110011101010: M1r = 2'b00;
			14'b00000111101010: M1r = 2'b00;
			14'b01000111101010: M1r = 2'b00;
			14'b10000111101010: M1r = 2'b01;
			14'b11000111101010: M1r = 2'b01;
			14'b00010111101010: M1r = 2'b00;
			14'b01010111101010: M1r = 2'b00;
			14'b10010111101010: M1r = 2'b00;
			14'b11010111101010: M1r = 2'b00;
			14'b00100111101010: M1r = 2'b00;
			14'b01100111101010: M1r = 2'b00;
			14'b10100111101010: M1r = 2'b00;
			14'b11100111101010: M1r = 2'b00;
			14'b00110111101010: M1r = 2'b00;
			14'b01110111101010: M1r = 2'b00;
			14'b10110111101010: M1r = 2'b00;
			14'b11110111101010: M1r = 2'b00;
			14'b00001011101010: M1r = 2'b01;
			14'b01001011101010: M1r = 2'b01;
			14'b10001011101010: M1r = 2'b01;
			14'b11001011101010: M1r = 2'b10;
			14'b00011011101010: M1r = 2'b01;
			14'b01011011101010: M1r = 2'b01;
			14'b10011011101010: M1r = 2'b01;
			14'b11011011101010: M1r = 2'b01;
			14'b00101011101010: M1r = 2'b00;
			14'b01101011101010: M1r = 2'b00;
			14'b10101011101010: M1r = 2'b00;
			14'b11101011101010: M1r = 2'b01;
			14'b00111011101010: M1r = 2'b00;
			14'b01111011101010: M1r = 2'b00;
			14'b10111011101010: M1r = 2'b00;
			14'b11111011101010: M1r = 2'b00;
			14'b00001111101010: M1r = 2'b10;
			14'b01001111101010: M1r = 2'b10;
			14'b10001111101010: M1r = 2'b10;
			14'b11001111101010: M1r = 2'b10;
			14'b00011111101010: M1r = 2'b01;
			14'b01011111101010: M1r = 2'b01;
			14'b10011111101010: M1r = 2'b10;
			14'b11011111101010: M1r = 2'b10;
			14'b00101111101010: M1r = 2'b01;
			14'b01101111101010: M1r = 2'b01;
			14'b10101111101010: M1r = 2'b01;
			14'b11101111101010: M1r = 2'b01;
			14'b00111111101010: M1r = 2'b00;
			14'b01111111101010: M1r = 2'b01;
			14'b10111111101010: M1r = 2'b01;
			14'b11111111101010: M1r = 2'b01;
			14'b00000000111010: M1r = 2'b01;
			14'b01000000111010: M1r = 2'b01;
			14'b10000000111010: M1r = 2'b01;
			14'b11000000111010: M1r = 2'b01;
			14'b00010000111010: M1r = 2'b00;
			14'b01010000111010: M1r = 2'b00;
			14'b10010000111010: M1r = 2'b01;
			14'b11010000111010: M1r = 2'b01;
			14'b00100000111010: M1r = 2'b00;
			14'b01100000111010: M1r = 2'b00;
			14'b10100000111010: M1r = 2'b00;
			14'b11100000111010: M1r = 2'b00;
			14'b00110000111010: M1r = 2'b00;
			14'b01110000111010: M1r = 2'b00;
			14'b10110000111010: M1r = 2'b00;
			14'b11110000111010: M1r = 2'b00;
			14'b00000100111010: M1r = 2'b10;
			14'b01000100111010: M1r = 2'b10;
			14'b10000100111010: M1r = 2'b10;
			14'b11000100111010: M1r = 2'b10;
			14'b00010100111010: M1r = 2'b01;
			14'b01010100111010: M1r = 2'b01;
			14'b10010100111010: M1r = 2'b01;
			14'b11010100111010: M1r = 2'b10;
			14'b00100100111010: M1r = 2'b01;
			14'b01100100111010: M1r = 2'b01;
			14'b10100100111010: M1r = 2'b01;
			14'b11100100111010: M1r = 2'b01;
			14'b00110100111010: M1r = 2'b00;
			14'b01110100111010: M1r = 2'b00;
			14'b10110100111010: M1r = 2'b00;
			14'b11110100111010: M1r = 2'b01;
			14'b00001000111010: M1r = 2'b10;
			14'b01001000111010: M1r = 2'b10;
			14'b10001000111010: M1r = 2'b11;
			14'b11001000111010: M1r = 2'b11;
			14'b00011000111010: M1r = 2'b10;
			14'b01011000111010: M1r = 2'b10;
			14'b10011000111010: M1r = 2'b10;
			14'b11011000111010: M1r = 2'b10;
			14'b00101000111010: M1r = 2'b01;
			14'b01101000111010: M1r = 2'b10;
			14'b10101000111010: M1r = 2'b10;
			14'b11101000111010: M1r = 2'b10;
			14'b00111000111010: M1r = 2'b01;
			14'b01111000111010: M1r = 2'b01;
			14'b10111000111010: M1r = 2'b01;
			14'b11111000111010: M1r = 2'b01;
			14'b00001100111010: M1r = 2'b11;
			14'b01001100111010: M1r = 2'b11;
			14'b10001100111010: M1r = 2'b11;
			14'b11001100111010: M1r = 2'b11;
			14'b00011100111010: M1r = 2'b11;
			14'b01011100111010: M1r = 2'b11;
			14'b10011100111010: M1r = 2'b11;
			14'b11011100111010: M1r = 2'b11;
			14'b00101100111010: M1r = 2'b10;
			14'b01101100111010: M1r = 2'b10;
			14'b10101100111010: M1r = 2'b10;
			14'b11101100111010: M1r = 2'b11;
			14'b00111100111010: M1r = 2'b10;
			14'b01111100111010: M1r = 2'b10;
			14'b10111100111010: M1r = 2'b10;
			14'b11111100111010: M1r = 2'b10;
			14'b00000001111010: M1r = 2'b01;
			14'b01000001111010: M1r = 2'b01;
			14'b10000001111010: M1r = 2'b01;
			14'b11000001111010: M1r = 2'b01;
			14'b00010001111010: M1r = 2'b00;
			14'b01010001111010: M1r = 2'b00;
			14'b10010001111010: M1r = 2'b00;
			14'b11010001111010: M1r = 2'b01;
			14'b00100001111010: M1r = 2'b00;
			14'b01100001111010: M1r = 2'b00;
			14'b10100001111010: M1r = 2'b00;
			14'b11100001111010: M1r = 2'b00;
			14'b00110001111010: M1r = 2'b00;
			14'b01110001111010: M1r = 2'b00;
			14'b10110001111010: M1r = 2'b00;
			14'b11110001111010: M1r = 2'b00;
			14'b00000101111010: M1r = 2'b01;
			14'b01000101111010: M1r = 2'b01;
			14'b10000101111010: M1r = 2'b10;
			14'b11000101111010: M1r = 2'b10;
			14'b00010101111010: M1r = 2'b01;
			14'b01010101111010: M1r = 2'b01;
			14'b10010101111010: M1r = 2'b01;
			14'b11010101111010: M1r = 2'b01;
			14'b00100101111010: M1r = 2'b00;
			14'b01100101111010: M1r = 2'b00;
			14'b10100101111010: M1r = 2'b01;
			14'b11100101111010: M1r = 2'b01;
			14'b00110101111010: M1r = 2'b00;
			14'b01110101111010: M1r = 2'b00;
			14'b10110101111010: M1r = 2'b00;
			14'b11110101111010: M1r = 2'b00;
			14'b00001001111010: M1r = 2'b10;
			14'b01001001111010: M1r = 2'b10;
			14'b10001001111010: M1r = 2'b10;
			14'b11001001111010: M1r = 2'b11;
			14'b00011001111010: M1r = 2'b10;
			14'b01011001111010: M1r = 2'b10;
			14'b10011001111010: M1r = 2'b10;
			14'b11011001111010: M1r = 2'b10;
			14'b00101001111010: M1r = 2'b01;
			14'b01101001111010: M1r = 2'b01;
			14'b10101001111010: M1r = 2'b01;
			14'b11101001111010: M1r = 2'b10;
			14'b00111001111010: M1r = 2'b01;
			14'b01111001111010: M1r = 2'b01;
			14'b10111001111010: M1r = 2'b01;
			14'b11111001111010: M1r = 2'b01;
			14'b00001101111010: M1r = 2'b11;
			14'b01001101111010: M1r = 2'b11;
			14'b10001101111010: M1r = 2'b11;
			14'b11001101111010: M1r = 2'b11;
			14'b00011101111010: M1r = 2'b10;
			14'b01011101111010: M1r = 2'b10;
			14'b10011101111010: M1r = 2'b11;
			14'b11011101111010: M1r = 2'b11;
			14'b00101101111010: M1r = 2'b10;
			14'b01101101111010: M1r = 2'b10;
			14'b10101101111010: M1r = 2'b10;
			14'b11101101111010: M1r = 2'b10;
			14'b00111101111010: M1r = 2'b01;
			14'b01111101111010: M1r = 2'b10;
			14'b10111101111010: M1r = 2'b10;
			14'b11111101111010: M1r = 2'b10;
			14'b00000010111010: M1r = 2'b00;
			14'b01000010111010: M1r = 2'b00;
			14'b10000010111010: M1r = 2'b01;
			14'b11000010111010: M1r = 2'b01;
			14'b00010010111010: M1r = 2'b00;
			14'b01010010111010: M1r = 2'b00;
			14'b10010010111010: M1r = 2'b00;
			14'b11010010111010: M1r = 2'b00;
			14'b00100010111010: M1r = 2'b00;
			14'b01100010111010: M1r = 2'b00;
			14'b10100010111010: M1r = 2'b00;
			14'b11100010111010: M1r = 2'b00;
			14'b00110010111010: M1r = 2'b00;
			14'b01110010111010: M1r = 2'b00;
			14'b10110010111010: M1r = 2'b00;
			14'b11110010111010: M1r = 2'b00;
			14'b00000110111010: M1r = 2'b01;
			14'b01000110111010: M1r = 2'b01;
			14'b10000110111010: M1r = 2'b01;
			14'b11000110111010: M1r = 2'b01;
			14'b00010110111010: M1r = 2'b01;
			14'b01010110111010: M1r = 2'b01;
			14'b10010110111010: M1r = 2'b01;
			14'b11010110111010: M1r = 2'b01;
			14'b00100110111010: M1r = 2'b00;
			14'b01100110111010: M1r = 2'b00;
			14'b10100110111010: M1r = 2'b00;
			14'b11100110111010: M1r = 2'b01;
			14'b00110110111010: M1r = 2'b00;
			14'b01110110111010: M1r = 2'b00;
			14'b10110110111010: M1r = 2'b00;
			14'b11110110111010: M1r = 2'b00;
			14'b00001010111010: M1r = 2'b10;
			14'b01001010111010: M1r = 2'b10;
			14'b10001010111010: M1r = 2'b10;
			14'b11001010111010: M1r = 2'b10;
			14'b00011010111010: M1r = 2'b01;
			14'b01011010111010: M1r = 2'b01;
			14'b10011010111010: M1r = 2'b10;
			14'b11011010111010: M1r = 2'b10;
			14'b00101010111010: M1r = 2'b01;
			14'b01101010111010: M1r = 2'b01;
			14'b10101010111010: M1r = 2'b01;
			14'b11101010111010: M1r = 2'b01;
			14'b00111010111010: M1r = 2'b00;
			14'b01111010111010: M1r = 2'b00;
			14'b10111010111010: M1r = 2'b01;
			14'b11111010111010: M1r = 2'b01;
			14'b00001110111010: M1r = 2'b11;
			14'b01001110111010: M1r = 2'b11;
			14'b10001110111010: M1r = 2'b11;
			14'b11001110111010: M1r = 2'b11;
			14'b00011110111010: M1r = 2'b10;
			14'b01011110111010: M1r = 2'b10;
			14'b10011110111010: M1r = 2'b10;
			14'b11011110111010: M1r = 2'b11;
			14'b00101110111010: M1r = 2'b10;
			14'b01101110111010: M1r = 2'b10;
			14'b10101110111010: M1r = 2'b10;
			14'b11101110111010: M1r = 2'b10;
			14'b00111110111010: M1r = 2'b01;
			14'b01111110111010: M1r = 2'b01;
			14'b10111110111010: M1r = 2'b01;
			14'b11111110111010: M1r = 2'b10;
			14'b00000011111010: M1r = 2'b00;
			14'b01000011111010: M1r = 2'b00;
			14'b10000011111010: M1r = 2'b00;
			14'b11000011111010: M1r = 2'b00;
			14'b00010011111010: M1r = 2'b00;
			14'b01010011111010: M1r = 2'b00;
			14'b10010011111010: M1r = 2'b00;
			14'b11010011111010: M1r = 2'b00;
			14'b00100011111010: M1r = 2'b00;
			14'b01100011111010: M1r = 2'b00;
			14'b10100011111010: M1r = 2'b00;
			14'b11100011111010: M1r = 2'b00;
			14'b00110011111010: M1r = 2'b00;
			14'b01110011111010: M1r = 2'b00;
			14'b10110011111010: M1r = 2'b00;
			14'b11110011111010: M1r = 2'b00;
			14'b00000111111010: M1r = 2'b01;
			14'b01000111111010: M1r = 2'b01;
			14'b10000111111010: M1r = 2'b01;
			14'b11000111111010: M1r = 2'b01;
			14'b00010111111010: M1r = 2'b00;
			14'b01010111111010: M1r = 2'b00;
			14'b10010111111010: M1r = 2'b01;
			14'b11010111111010: M1r = 2'b01;
			14'b00100111111010: M1r = 2'b00;
			14'b01100111111010: M1r = 2'b00;
			14'b10100111111010: M1r = 2'b00;
			14'b11100111111010: M1r = 2'b00;
			14'b00110111111010: M1r = 2'b00;
			14'b01110111111010: M1r = 2'b00;
			14'b10110111111010: M1r = 2'b00;
			14'b11110111111010: M1r = 2'b00;
			14'b00001011111010: M1r = 2'b01;
			14'b01001011111010: M1r = 2'b10;
			14'b10001011111010: M1r = 2'b10;
			14'b11001011111010: M1r = 2'b10;
			14'b00011011111010: M1r = 2'b01;
			14'b01011011111010: M1r = 2'b01;
			14'b10011011111010: M1r = 2'b01;
			14'b11011011111010: M1r = 2'b01;
			14'b00101011111010: M1r = 2'b01;
			14'b01101011111010: M1r = 2'b01;
			14'b10101011111010: M1r = 2'b01;
			14'b11101011111010: M1r = 2'b01;
			14'b00111011111010: M1r = 2'b00;
			14'b01111011111010: M1r = 2'b00;
			14'b10111011111010: M1r = 2'b00;
			14'b11111011111010: M1r = 2'b01;
			14'b00001111111010: M1r = 2'b10;
			14'b01001111111010: M1r = 2'b10;
			14'b10001111111010: M1r = 2'b11;
			14'b11001111111010: M1r = 2'b11;
			14'b00011111111010: M1r = 2'b10;
			14'b01011111111010: M1r = 2'b10;
			14'b10011111111010: M1r = 2'b10;
			14'b11011111111010: M1r = 2'b10;
			14'b00101111111010: M1r = 2'b01;
			14'b01101111111010: M1r = 2'b01;
			14'b10101111111010: M1r = 2'b10;
			14'b11101111111010: M1r = 2'b10;
			14'b00111111111010: M1r = 2'b01;
			14'b01111111111010: M1r = 2'b01;
			14'b10111111111010: M1r = 2'b01;
			14'b11111111111010: M1r = 2'b01;
			14'b00000000001110: M1r = 2'b00;
			14'b01000000001110: M1r = 2'b00;
			14'b10000000001110: M1r = 2'b00;
			14'b11000000001110: M1r = 2'b00;
			14'b00010000001110: M1r = 2'b00;
			14'b01010000001110: M1r = 2'b00;
			14'b10010000001110: M1r = 2'b00;
			14'b11010000001110: M1r = 2'b00;
			14'b00100000001110: M1r = 2'b00;
			14'b01100000001110: M1r = 2'b00;
			14'b10100000001110: M1r = 2'b00;
			14'b11100000001110: M1r = 2'b00;
			14'b00110000001110: M1r = 2'b00;
			14'b01110000001110: M1r = 2'b00;
			14'b10110000001110: M1r = 2'b00;
			14'b11110000001110: M1r = 2'b00;
			14'b00000100001110: M1r = 2'b00;
			14'b01000100001110: M1r = 2'b00;
			14'b10000100001110: M1r = 2'b00;
			14'b11000100001110: M1r = 2'b00;
			14'b00010100001110: M1r = 2'b00;
			14'b01010100001110: M1r = 2'b00;
			14'b10010100001110: M1r = 2'b00;
			14'b11010100001110: M1r = 2'b00;
			14'b00100100001110: M1r = 2'b00;
			14'b01100100001110: M1r = 2'b00;
			14'b10100100001110: M1r = 2'b00;
			14'b11100100001110: M1r = 2'b00;
			14'b00110100001110: M1r = 2'b00;
			14'b01110100001110: M1r = 2'b00;
			14'b10110100001110: M1r = 2'b00;
			14'b11110100001110: M1r = 2'b00;
			14'b00001000001110: M1r = 2'b00;
			14'b01001000001110: M1r = 2'b00;
			14'b10001000001110: M1r = 2'b01;
			14'b11001000001110: M1r = 2'b01;
			14'b00011000001110: M1r = 2'b00;
			14'b01011000001110: M1r = 2'b00;
			14'b10011000001110: M1r = 2'b00;
			14'b11011000001110: M1r = 2'b00;
			14'b00101000001110: M1r = 2'b00;
			14'b01101000001110: M1r = 2'b00;
			14'b10101000001110: M1r = 2'b00;
			14'b11101000001110: M1r = 2'b00;
			14'b00111000001110: M1r = 2'b00;
			14'b01111000001110: M1r = 2'b00;
			14'b10111000001110: M1r = 2'b00;
			14'b11111000001110: M1r = 2'b00;
			14'b00001100001110: M1r = 2'b01;
			14'b01001100001110: M1r = 2'b01;
			14'b10001100001110: M1r = 2'b01;
			14'b11001100001110: M1r = 2'b01;
			14'b00011100001110: M1r = 2'b01;
			14'b01011100001110: M1r = 2'b01;
			14'b10011100001110: M1r = 2'b01;
			14'b11011100001110: M1r = 2'b01;
			14'b00101100001110: M1r = 2'b00;
			14'b01101100001110: M1r = 2'b00;
			14'b10101100001110: M1r = 2'b00;
			14'b11101100001110: M1r = 2'b01;
			14'b00111100001110: M1r = 2'b00;
			14'b01111100001110: M1r = 2'b00;
			14'b10111100001110: M1r = 2'b00;
			14'b11111100001110: M1r = 2'b00;
			14'b00000001001110: M1r = 2'b00;
			14'b01000001001110: M1r = 2'b00;
			14'b10000001001110: M1r = 2'b00;
			14'b11000001001110: M1r = 2'b00;
			14'b00010001001110: M1r = 2'b00;
			14'b01010001001110: M1r = 2'b00;
			14'b10010001001110: M1r = 2'b00;
			14'b11010001001110: M1r = 2'b00;
			14'b00100001001110: M1r = 2'b00;
			14'b01100001001110: M1r = 2'b00;
			14'b10100001001110: M1r = 2'b00;
			14'b11100001001110: M1r = 2'b00;
			14'b00110001001110: M1r = 2'b00;
			14'b01110001001110: M1r = 2'b00;
			14'b10110001001110: M1r = 2'b00;
			14'b11110001001110: M1r = 2'b00;
			14'b00000101001110: M1r = 2'b00;
			14'b01000101001110: M1r = 2'b00;
			14'b10000101001110: M1r = 2'b00;
			14'b11000101001110: M1r = 2'b00;
			14'b00010101001110: M1r = 2'b00;
			14'b01010101001110: M1r = 2'b00;
			14'b10010101001110: M1r = 2'b00;
			14'b11010101001110: M1r = 2'b00;
			14'b00100101001110: M1r = 2'b00;
			14'b01100101001110: M1r = 2'b00;
			14'b10100101001110: M1r = 2'b00;
			14'b11100101001110: M1r = 2'b00;
			14'b00110101001110: M1r = 2'b00;
			14'b01110101001110: M1r = 2'b00;
			14'b10110101001110: M1r = 2'b00;
			14'b11110101001110: M1r = 2'b00;
			14'b00001001001110: M1r = 2'b00;
			14'b01001001001110: M1r = 2'b00;
			14'b10001001001110: M1r = 2'b00;
			14'b11001001001110: M1r = 2'b00;
			14'b00011001001110: M1r = 2'b00;
			14'b01011001001110: M1r = 2'b00;
			14'b10011001001110: M1r = 2'b00;
			14'b11011001001110: M1r = 2'b00;
			14'b00101001001110: M1r = 2'b00;
			14'b01101001001110: M1r = 2'b00;
			14'b10101001001110: M1r = 2'b00;
			14'b11101001001110: M1r = 2'b00;
			14'b00111001001110: M1r = 2'b00;
			14'b01111001001110: M1r = 2'b00;
			14'b10111001001110: M1r = 2'b00;
			14'b11111001001110: M1r = 2'b00;
			14'b00001101001110: M1r = 2'b01;
			14'b01001101001110: M1r = 2'b01;
			14'b10001101001110: M1r = 2'b01;
			14'b11001101001110: M1r = 2'b01;
			14'b00011101001110: M1r = 2'b00;
			14'b01011101001110: M1r = 2'b00;
			14'b10011101001110: M1r = 2'b01;
			14'b11011101001110: M1r = 2'b01;
			14'b00101101001110: M1r = 2'b00;
			14'b01101101001110: M1r = 2'b00;
			14'b10101101001110: M1r = 2'b00;
			14'b11101101001110: M1r = 2'b00;
			14'b00111101001110: M1r = 2'b00;
			14'b01111101001110: M1r = 2'b00;
			14'b10111101001110: M1r = 2'b00;
			14'b11111101001110: M1r = 2'b00;
			14'b00000010001110: M1r = 2'b00;
			14'b01000010001110: M1r = 2'b00;
			14'b10000010001110: M1r = 2'b00;
			14'b11000010001110: M1r = 2'b00;
			14'b00010010001110: M1r = 2'b00;
			14'b01010010001110: M1r = 2'b00;
			14'b10010010001110: M1r = 2'b00;
			14'b11010010001110: M1r = 2'b00;
			14'b00100010001110: M1r = 2'b00;
			14'b01100010001110: M1r = 2'b00;
			14'b10100010001110: M1r = 2'b00;
			14'b11100010001110: M1r = 2'b00;
			14'b00110010001110: M1r = 2'b00;
			14'b01110010001110: M1r = 2'b00;
			14'b10110010001110: M1r = 2'b00;
			14'b11110010001110: M1r = 2'b00;
			14'b00000110001110: M1r = 2'b00;
			14'b01000110001110: M1r = 2'b00;
			14'b10000110001110: M1r = 2'b00;
			14'b11000110001110: M1r = 2'b00;
			14'b00010110001110: M1r = 2'b00;
			14'b01010110001110: M1r = 2'b00;
			14'b10010110001110: M1r = 2'b00;
			14'b11010110001110: M1r = 2'b00;
			14'b00100110001110: M1r = 2'b00;
			14'b01100110001110: M1r = 2'b00;
			14'b10100110001110: M1r = 2'b00;
			14'b11100110001110: M1r = 2'b00;
			14'b00110110001110: M1r = 2'b00;
			14'b01110110001110: M1r = 2'b00;
			14'b10110110001110: M1r = 2'b00;
			14'b11110110001110: M1r = 2'b00;
			14'b00001010001110: M1r = 2'b00;
			14'b01001010001110: M1r = 2'b00;
			14'b10001010001110: M1r = 2'b00;
			14'b11001010001110: M1r = 2'b00;
			14'b00011010001110: M1r = 2'b00;
			14'b01011010001110: M1r = 2'b00;
			14'b10011010001110: M1r = 2'b00;
			14'b11011010001110: M1r = 2'b00;
			14'b00101010001110: M1r = 2'b00;
			14'b01101010001110: M1r = 2'b00;
			14'b10101010001110: M1r = 2'b00;
			14'b11101010001110: M1r = 2'b00;
			14'b00111010001110: M1r = 2'b00;
			14'b01111010001110: M1r = 2'b00;
			14'b10111010001110: M1r = 2'b00;
			14'b11111010001110: M1r = 2'b00;
			14'b00001110001110: M1r = 2'b00;
			14'b01001110001110: M1r = 2'b01;
			14'b10001110001110: M1r = 2'b01;
			14'b11001110001110: M1r = 2'b01;
			14'b00011110001110: M1r = 2'b00;
			14'b01011110001110: M1r = 2'b00;
			14'b10011110001110: M1r = 2'b00;
			14'b11011110001110: M1r = 2'b00;
			14'b00101110001110: M1r = 2'b00;
			14'b01101110001110: M1r = 2'b00;
			14'b10101110001110: M1r = 2'b00;
			14'b11101110001110: M1r = 2'b00;
			14'b00111110001110: M1r = 2'b00;
			14'b01111110001110: M1r = 2'b00;
			14'b10111110001110: M1r = 2'b00;
			14'b11111110001110: M1r = 2'b00;
			14'b00000011001110: M1r = 2'b00;
			14'b01000011001110: M1r = 2'b00;
			14'b10000011001110: M1r = 2'b00;
			14'b11000011001110: M1r = 2'b00;
			14'b00010011001110: M1r = 2'b00;
			14'b01010011001110: M1r = 2'b00;
			14'b10010011001110: M1r = 2'b00;
			14'b11010011001110: M1r = 2'b00;
			14'b00100011001110: M1r = 2'b00;
			14'b01100011001110: M1r = 2'b00;
			14'b10100011001110: M1r = 2'b00;
			14'b11100011001110: M1r = 2'b00;
			14'b00110011001110: M1r = 2'b00;
			14'b01110011001110: M1r = 2'b00;
			14'b10110011001110: M1r = 2'b00;
			14'b11110011001110: M1r = 2'b00;
			14'b00000111001110: M1r = 2'b00;
			14'b01000111001110: M1r = 2'b00;
			14'b10000111001110: M1r = 2'b00;
			14'b11000111001110: M1r = 2'b00;
			14'b00010111001110: M1r = 2'b00;
			14'b01010111001110: M1r = 2'b00;
			14'b10010111001110: M1r = 2'b00;
			14'b11010111001110: M1r = 2'b00;
			14'b00100111001110: M1r = 2'b00;
			14'b01100111001110: M1r = 2'b00;
			14'b10100111001110: M1r = 2'b00;
			14'b11100111001110: M1r = 2'b00;
			14'b00110111001110: M1r = 2'b00;
			14'b01110111001110: M1r = 2'b00;
			14'b10110111001110: M1r = 2'b00;
			14'b11110111001110: M1r = 2'b00;
			14'b00001011001110: M1r = 2'b00;
			14'b01001011001110: M1r = 2'b00;
			14'b10001011001110: M1r = 2'b00;
			14'b11001011001110: M1r = 2'b00;
			14'b00011011001110: M1r = 2'b00;
			14'b01011011001110: M1r = 2'b00;
			14'b10011011001110: M1r = 2'b00;
			14'b11011011001110: M1r = 2'b00;
			14'b00101011001110: M1r = 2'b00;
			14'b01101011001110: M1r = 2'b00;
			14'b10101011001110: M1r = 2'b00;
			14'b11101011001110: M1r = 2'b00;
			14'b00111011001110: M1r = 2'b00;
			14'b01111011001110: M1r = 2'b00;
			14'b10111011001110: M1r = 2'b00;
			14'b11111011001110: M1r = 2'b00;
			14'b00001111001110: M1r = 2'b00;
			14'b01001111001110: M1r = 2'b00;
			14'b10001111001110: M1r = 2'b00;
			14'b11001111001110: M1r = 2'b01;
			14'b00011111001110: M1r = 2'b00;
			14'b01011111001110: M1r = 2'b00;
			14'b10011111001110: M1r = 2'b00;
			14'b11011111001110: M1r = 2'b00;
			14'b00101111001110: M1r = 2'b00;
			14'b01101111001110: M1r = 2'b00;
			14'b10101111001110: M1r = 2'b00;
			14'b11101111001110: M1r = 2'b00;
			14'b00111111001110: M1r = 2'b00;
			14'b01111111001110: M1r = 2'b00;
			14'b10111111001110: M1r = 2'b00;
			14'b11111111001110: M1r = 2'b00;
			14'b00000000011110: M1r = 2'b00;
			14'b01000000011110: M1r = 2'b00;
			14'b10000000011110: M1r = 2'b00;
			14'b11000000011110: M1r = 2'b00;
			14'b00010000011110: M1r = 2'b00;
			14'b01010000011110: M1r = 2'b00;
			14'b10010000011110: M1r = 2'b00;
			14'b11010000011110: M1r = 2'b00;
			14'b00100000011110: M1r = 2'b00;
			14'b01100000011110: M1r = 2'b00;
			14'b10100000011110: M1r = 2'b00;
			14'b11100000011110: M1r = 2'b00;
			14'b00110000011110: M1r = 2'b00;
			14'b01110000011110: M1r = 2'b00;
			14'b10110000011110: M1r = 2'b00;
			14'b11110000011110: M1r = 2'b00;
			14'b00000100011110: M1r = 2'b00;
			14'b01000100011110: M1r = 2'b00;
			14'b10000100011110: M1r = 2'b00;
			14'b11000100011110: M1r = 2'b00;
			14'b00010100011110: M1r = 2'b00;
			14'b01010100011110: M1r = 2'b00;
			14'b10010100011110: M1r = 2'b00;
			14'b11010100011110: M1r = 2'b00;
			14'b00100100011110: M1r = 2'b00;
			14'b01100100011110: M1r = 2'b00;
			14'b10100100011110: M1r = 2'b00;
			14'b11100100011110: M1r = 2'b00;
			14'b00110100011110: M1r = 2'b00;
			14'b01110100011110: M1r = 2'b00;
			14'b10110100011110: M1r = 2'b00;
			14'b11110100011110: M1r = 2'b00;
			14'b00001000011110: M1r = 2'b01;
			14'b01001000011110: M1r = 2'b01;
			14'b10001000011110: M1r = 2'b01;
			14'b11001000011110: M1r = 2'b01;
			14'b00011000011110: M1r = 2'b00;
			14'b01011000011110: M1r = 2'b00;
			14'b10011000011110: M1r = 2'b01;
			14'b11011000011110: M1r = 2'b01;
			14'b00101000011110: M1r = 2'b00;
			14'b01101000011110: M1r = 2'b00;
			14'b10101000011110: M1r = 2'b00;
			14'b11101000011110: M1r = 2'b00;
			14'b00111000011110: M1r = 2'b00;
			14'b01111000011110: M1r = 2'b00;
			14'b10111000011110: M1r = 2'b00;
			14'b11111000011110: M1r = 2'b00;
			14'b00001100011110: M1r = 2'b01;
			14'b01001100011110: M1r = 2'b10;
			14'b10001100011110: M1r = 2'b10;
			14'b11001100011110: M1r = 2'b10;
			14'b00011100011110: M1r = 2'b01;
			14'b01011100011110: M1r = 2'b01;
			14'b10011100011110: M1r = 2'b01;
			14'b11011100011110: M1r = 2'b01;
			14'b00101100011110: M1r = 2'b00;
			14'b01101100011110: M1r = 2'b01;
			14'b10101100011110: M1r = 2'b01;
			14'b11101100011110: M1r = 2'b01;
			14'b00111100011110: M1r = 2'b00;
			14'b01111100011110: M1r = 2'b00;
			14'b10111100011110: M1r = 2'b00;
			14'b11111100011110: M1r = 2'b00;
			14'b00000001011110: M1r = 2'b00;
			14'b01000001011110: M1r = 2'b00;
			14'b10000001011110: M1r = 2'b00;
			14'b11000001011110: M1r = 2'b00;
			14'b00010001011110: M1r = 2'b00;
			14'b01010001011110: M1r = 2'b00;
			14'b10010001011110: M1r = 2'b00;
			14'b11010001011110: M1r = 2'b00;
			14'b00100001011110: M1r = 2'b00;
			14'b01100001011110: M1r = 2'b00;
			14'b10100001011110: M1r = 2'b00;
			14'b11100001011110: M1r = 2'b00;
			14'b00110001011110: M1r = 2'b00;
			14'b01110001011110: M1r = 2'b00;
			14'b10110001011110: M1r = 2'b00;
			14'b11110001011110: M1r = 2'b00;
			14'b00000101011110: M1r = 2'b00;
			14'b01000101011110: M1r = 2'b00;
			14'b10000101011110: M1r = 2'b00;
			14'b11000101011110: M1r = 2'b00;
			14'b00010101011110: M1r = 2'b00;
			14'b01010101011110: M1r = 2'b00;
			14'b10010101011110: M1r = 2'b00;
			14'b11010101011110: M1r = 2'b00;
			14'b00100101011110: M1r = 2'b00;
			14'b01100101011110: M1r = 2'b00;
			14'b10100101011110: M1r = 2'b00;
			14'b11100101011110: M1r = 2'b00;
			14'b00110101011110: M1r = 2'b00;
			14'b01110101011110: M1r = 2'b00;
			14'b10110101011110: M1r = 2'b00;
			14'b11110101011110: M1r = 2'b00;
			14'b00001001011110: M1r = 2'b00;
			14'b01001001011110: M1r = 2'b01;
			14'b10001001011110: M1r = 2'b01;
			14'b11001001011110: M1r = 2'b01;
			14'b00011001011110: M1r = 2'b00;
			14'b01011001011110: M1r = 2'b00;
			14'b10011001011110: M1r = 2'b00;
			14'b11011001011110: M1r = 2'b00;
			14'b00101001011110: M1r = 2'b00;
			14'b01101001011110: M1r = 2'b00;
			14'b10101001011110: M1r = 2'b00;
			14'b11101001011110: M1r = 2'b00;
			14'b00111001011110: M1r = 2'b00;
			14'b01111001011110: M1r = 2'b00;
			14'b10111001011110: M1r = 2'b00;
			14'b11111001011110: M1r = 2'b00;
			14'b00001101011110: M1r = 2'b01;
			14'b01001101011110: M1r = 2'b01;
			14'b10001101011110: M1r = 2'b01;
			14'b11001101011110: M1r = 2'b10;
			14'b00011101011110: M1r = 2'b01;
			14'b01011101011110: M1r = 2'b01;
			14'b10011101011110: M1r = 2'b01;
			14'b11011101011110: M1r = 2'b01;
			14'b00101101011110: M1r = 2'b00;
			14'b01101101011110: M1r = 2'b00;
			14'b10101101011110: M1r = 2'b01;
			14'b11101101011110: M1r = 2'b01;
			14'b00111101011110: M1r = 2'b00;
			14'b01111101011110: M1r = 2'b00;
			14'b10111101011110: M1r = 2'b00;
			14'b11111101011110: M1r = 2'b00;
			14'b00000010011110: M1r = 2'b00;
			14'b01000010011110: M1r = 2'b00;
			14'b10000010011110: M1r = 2'b00;
			14'b11000010011110: M1r = 2'b00;
			14'b00010010011110: M1r = 2'b00;
			14'b01010010011110: M1r = 2'b00;
			14'b10010010011110: M1r = 2'b00;
			14'b11010010011110: M1r = 2'b00;
			14'b00100010011110: M1r = 2'b00;
			14'b01100010011110: M1r = 2'b00;
			14'b10100010011110: M1r = 2'b00;
			14'b11100010011110: M1r = 2'b00;
			14'b00110010011110: M1r = 2'b00;
			14'b01110010011110: M1r = 2'b00;
			14'b10110010011110: M1r = 2'b00;
			14'b11110010011110: M1r = 2'b00;
			14'b00000110011110: M1r = 2'b00;
			14'b01000110011110: M1r = 2'b00;
			14'b10000110011110: M1r = 2'b00;
			14'b11000110011110: M1r = 2'b00;
			14'b00010110011110: M1r = 2'b00;
			14'b01010110011110: M1r = 2'b00;
			14'b10010110011110: M1r = 2'b00;
			14'b11010110011110: M1r = 2'b00;
			14'b00100110011110: M1r = 2'b00;
			14'b01100110011110: M1r = 2'b00;
			14'b10100110011110: M1r = 2'b00;
			14'b11100110011110: M1r = 2'b00;
			14'b00110110011110: M1r = 2'b00;
			14'b01110110011110: M1r = 2'b00;
			14'b10110110011110: M1r = 2'b00;
			14'b11110110011110: M1r = 2'b00;
			14'b00001010011110: M1r = 2'b00;
			14'b01001010011110: M1r = 2'b00;
			14'b10001010011110: M1r = 2'b00;
			14'b11001010011110: M1r = 2'b01;
			14'b00011010011110: M1r = 2'b00;
			14'b01011010011110: M1r = 2'b00;
			14'b10011010011110: M1r = 2'b00;
			14'b11011010011110: M1r = 2'b00;
			14'b00101010011110: M1r = 2'b00;
			14'b01101010011110: M1r = 2'b00;
			14'b10101010011110: M1r = 2'b00;
			14'b11101010011110: M1r = 2'b00;
			14'b00111010011110: M1r = 2'b00;
			14'b01111010011110: M1r = 2'b00;
			14'b10111010011110: M1r = 2'b00;
			14'b11111010011110: M1r = 2'b00;
			14'b00001110011110: M1r = 2'b01;
			14'b01001110011110: M1r = 2'b01;
			14'b10001110011110: M1r = 2'b01;
			14'b11001110011110: M1r = 2'b01;
			14'b00011110011110: M1r = 2'b00;
			14'b01011110011110: M1r = 2'b01;
			14'b10011110011110: M1r = 2'b01;
			14'b11011110011110: M1r = 2'b01;
			14'b00101110011110: M1r = 2'b00;
			14'b01101110011110: M1r = 2'b00;
			14'b10101110011110: M1r = 2'b00;
			14'b11101110011110: M1r = 2'b00;
			14'b00111110011110: M1r = 2'b00;
			14'b01111110011110: M1r = 2'b00;
			14'b10111110011110: M1r = 2'b00;
			14'b11111110011110: M1r = 2'b00;
			14'b00000011011110: M1r = 2'b00;
			14'b01000011011110: M1r = 2'b00;
			14'b10000011011110: M1r = 2'b00;
			14'b11000011011110: M1r = 2'b00;
			14'b00010011011110: M1r = 2'b00;
			14'b01010011011110: M1r = 2'b00;
			14'b10010011011110: M1r = 2'b00;
			14'b11010011011110: M1r = 2'b00;
			14'b00100011011110: M1r = 2'b00;
			14'b01100011011110: M1r = 2'b00;
			14'b10100011011110: M1r = 2'b00;
			14'b11100011011110: M1r = 2'b00;
			14'b00110011011110: M1r = 2'b00;
			14'b01110011011110: M1r = 2'b00;
			14'b10110011011110: M1r = 2'b00;
			14'b11110011011110: M1r = 2'b00;
			14'b00000111011110: M1r = 2'b00;
			14'b01000111011110: M1r = 2'b00;
			14'b10000111011110: M1r = 2'b00;
			14'b11000111011110: M1r = 2'b00;
			14'b00010111011110: M1r = 2'b00;
			14'b01010111011110: M1r = 2'b00;
			14'b10010111011110: M1r = 2'b00;
			14'b11010111011110: M1r = 2'b00;
			14'b00100111011110: M1r = 2'b00;
			14'b01100111011110: M1r = 2'b00;
			14'b10100111011110: M1r = 2'b00;
			14'b11100111011110: M1r = 2'b00;
			14'b00110111011110: M1r = 2'b00;
			14'b01110111011110: M1r = 2'b00;
			14'b10110111011110: M1r = 2'b00;
			14'b11110111011110: M1r = 2'b00;
			14'b00001011011110: M1r = 2'b00;
			14'b01001011011110: M1r = 2'b00;
			14'b10001011011110: M1r = 2'b00;
			14'b11001011011110: M1r = 2'b00;
			14'b00011011011110: M1r = 2'b00;
			14'b01011011011110: M1r = 2'b00;
			14'b10011011011110: M1r = 2'b00;
			14'b11011011011110: M1r = 2'b00;
			14'b00101011011110: M1r = 2'b00;
			14'b01101011011110: M1r = 2'b00;
			14'b10101011011110: M1r = 2'b00;
			14'b11101011011110: M1r = 2'b00;
			14'b00111011011110: M1r = 2'b00;
			14'b01111011011110: M1r = 2'b00;
			14'b10111011011110: M1r = 2'b00;
			14'b11111011011110: M1r = 2'b00;
			14'b00001111011110: M1r = 2'b01;
			14'b01001111011110: M1r = 2'b01;
			14'b10001111011110: M1r = 2'b01;
			14'b11001111011110: M1r = 2'b01;
			14'b00011111011110: M1r = 2'b00;
			14'b01011111011110: M1r = 2'b00;
			14'b10011111011110: M1r = 2'b00;
			14'b11011111011110: M1r = 2'b01;
			14'b00101111011110: M1r = 2'b00;
			14'b01101111011110: M1r = 2'b00;
			14'b10101111011110: M1r = 2'b00;
			14'b11101111011110: M1r = 2'b00;
			14'b00111111011110: M1r = 2'b00;
			14'b01111111011110: M1r = 2'b00;
			14'b10111111011110: M1r = 2'b00;
			14'b11111111011110: M1r = 2'b00;
			14'b00000000101110: M1r = 2'b00;
			14'b01000000101110: M1r = 2'b00;
			14'b10000000101110: M1r = 2'b00;
			14'b11000000101110: M1r = 2'b00;
			14'b00010000101110: M1r = 2'b00;
			14'b01010000101110: M1r = 2'b00;
			14'b10010000101110: M1r = 2'b00;
			14'b11010000101110: M1r = 2'b00;
			14'b00100000101110: M1r = 2'b00;
			14'b01100000101110: M1r = 2'b00;
			14'b10100000101110: M1r = 2'b00;
			14'b11100000101110: M1r = 2'b00;
			14'b00110000101110: M1r = 2'b00;
			14'b01110000101110: M1r = 2'b00;
			14'b10110000101110: M1r = 2'b00;
			14'b11110000101110: M1r = 2'b00;
			14'b00000100101110: M1r = 2'b00;
			14'b01000100101110: M1r = 2'b01;
			14'b10000100101110: M1r = 2'b01;
			14'b11000100101110: M1r = 2'b01;
			14'b00010100101110: M1r = 2'b00;
			14'b01010100101110: M1r = 2'b00;
			14'b10010100101110: M1r = 2'b00;
			14'b11010100101110: M1r = 2'b00;
			14'b00100100101110: M1r = 2'b00;
			14'b01100100101110: M1r = 2'b00;
			14'b10100100101110: M1r = 2'b00;
			14'b11100100101110: M1r = 2'b00;
			14'b00110100101110: M1r = 2'b00;
			14'b01110100101110: M1r = 2'b00;
			14'b10110100101110: M1r = 2'b00;
			14'b11110100101110: M1r = 2'b00;
			14'b00001000101110: M1r = 2'b01;
			14'b01001000101110: M1r = 2'b01;
			14'b10001000101110: M1r = 2'b01;
			14'b11001000101110: M1r = 2'b10;
			14'b00011000101110: M1r = 2'b01;
			14'b01011000101110: M1r = 2'b01;
			14'b10011000101110: M1r = 2'b01;
			14'b11011000101110: M1r = 2'b01;
			14'b00101000101110: M1r = 2'b00;
			14'b01101000101110: M1r = 2'b00;
			14'b10101000101110: M1r = 2'b00;
			14'b11101000101110: M1r = 2'b01;
			14'b00111000101110: M1r = 2'b00;
			14'b01111000101110: M1r = 2'b00;
			14'b10111000101110: M1r = 2'b00;
			14'b11111000101110: M1r = 2'b00;
			14'b00001100101110: M1r = 2'b10;
			14'b01001100101110: M1r = 2'b10;
			14'b10001100101110: M1r = 2'b10;
			14'b11001100101110: M1r = 2'b10;
			14'b00011100101110: M1r = 2'b01;
			14'b01011100101110: M1r = 2'b10;
			14'b10011100101110: M1r = 2'b10;
			14'b11011100101110: M1r = 2'b10;
			14'b00101100101110: M1r = 2'b01;
			14'b01101100101110: M1r = 2'b01;
			14'b10101100101110: M1r = 2'b01;
			14'b11101100101110: M1r = 2'b01;
			14'b00111100101110: M1r = 2'b00;
			14'b01111100101110: M1r = 2'b01;
			14'b10111100101110: M1r = 2'b01;
			14'b11111100101110: M1r = 2'b01;
			14'b00000001101110: M1r = 2'b00;
			14'b01000001101110: M1r = 2'b00;
			14'b10000001101110: M1r = 2'b00;
			14'b11000001101110: M1r = 2'b00;
			14'b00010001101110: M1r = 2'b00;
			14'b01010001101110: M1r = 2'b00;
			14'b10010001101110: M1r = 2'b00;
			14'b11010001101110: M1r = 2'b00;
			14'b00100001101110: M1r = 2'b00;
			14'b01100001101110: M1r = 2'b00;
			14'b10100001101110: M1r = 2'b00;
			14'b11100001101110: M1r = 2'b00;
			14'b00110001101110: M1r = 2'b00;
			14'b01110001101110: M1r = 2'b00;
			14'b10110001101110: M1r = 2'b00;
			14'b11110001101110: M1r = 2'b00;
			14'b00000101101110: M1r = 2'b00;
			14'b01000101101110: M1r = 2'b00;
			14'b10000101101110: M1r = 2'b00;
			14'b11000101101110: M1r = 2'b01;
			14'b00010101101110: M1r = 2'b00;
			14'b01010101101110: M1r = 2'b00;
			14'b10010101101110: M1r = 2'b00;
			14'b11010101101110: M1r = 2'b00;
			14'b00100101101110: M1r = 2'b00;
			14'b01100101101110: M1r = 2'b00;
			14'b10100101101110: M1r = 2'b00;
			14'b11100101101110: M1r = 2'b00;
			14'b00110101101110: M1r = 2'b00;
			14'b01110101101110: M1r = 2'b00;
			14'b10110101101110: M1r = 2'b00;
			14'b11110101101110: M1r = 2'b00;
			14'b00001001101110: M1r = 2'b01;
			14'b01001001101110: M1r = 2'b01;
			14'b10001001101110: M1r = 2'b01;
			14'b11001001101110: M1r = 2'b01;
			14'b00011001101110: M1r = 2'b00;
			14'b01011001101110: M1r = 2'b01;
			14'b10011001101110: M1r = 2'b01;
			14'b11011001101110: M1r = 2'b01;
			14'b00101001101110: M1r = 2'b00;
			14'b01101001101110: M1r = 2'b00;
			14'b10101001101110: M1r = 2'b00;
			14'b11101001101110: M1r = 2'b00;
			14'b00111001101110: M1r = 2'b00;
			14'b01111001101110: M1r = 2'b00;
			14'b10111001101110: M1r = 2'b00;
			14'b11111001101110: M1r = 2'b00;
			14'b00001101101110: M1r = 2'b10;
			14'b01001101101110: M1r = 2'b10;
			14'b10001101101110: M1r = 2'b10;
			14'b11001101101110: M1r = 2'b10;
			14'b00011101101110: M1r = 2'b01;
			14'b01011101101110: M1r = 2'b01;
			14'b10011101101110: M1r = 2'b01;
			14'b11011101101110: M1r = 2'b10;
			14'b00101101101110: M1r = 2'b01;
			14'b01101101101110: M1r = 2'b01;
			14'b10101101101110: M1r = 2'b01;
			14'b11101101101110: M1r = 2'b01;
			14'b00111101101110: M1r = 2'b00;
			14'b01111101101110: M1r = 2'b00;
			14'b10111101101110: M1r = 2'b00;
			14'b11111101101110: M1r = 2'b01;
			14'b00000010101110: M1r = 2'b00;
			14'b01000010101110: M1r = 2'b00;
			14'b10000010101110: M1r = 2'b00;
			14'b11000010101110: M1r = 2'b00;
			14'b00010010101110: M1r = 2'b00;
			14'b01010010101110: M1r = 2'b00;
			14'b10010010101110: M1r = 2'b00;
			14'b11010010101110: M1r = 2'b00;
			14'b00100010101110: M1r = 2'b00;
			14'b01100010101110: M1r = 2'b00;
			14'b10100010101110: M1r = 2'b00;
			14'b11100010101110: M1r = 2'b00;
			14'b00110010101110: M1r = 2'b00;
			14'b01110010101110: M1r = 2'b00;
			14'b10110010101110: M1r = 2'b00;
			14'b11110010101110: M1r = 2'b00;
			14'b00000110101110: M1r = 2'b00;
			14'b01000110101110: M1r = 2'b00;
			14'b10000110101110: M1r = 2'b00;
			14'b11000110101110: M1r = 2'b00;
			14'b00010110101110: M1r = 2'b00;
			14'b01010110101110: M1r = 2'b00;
			14'b10010110101110: M1r = 2'b00;
			14'b11010110101110: M1r = 2'b00;
			14'b00100110101110: M1r = 2'b00;
			14'b01100110101110: M1r = 2'b00;
			14'b10100110101110: M1r = 2'b00;
			14'b11100110101110: M1r = 2'b00;
			14'b00110110101110: M1r = 2'b00;
			14'b01110110101110: M1r = 2'b00;
			14'b10110110101110: M1r = 2'b00;
			14'b11110110101110: M1r = 2'b00;
			14'b00001010101110: M1r = 2'b01;
			14'b01001010101110: M1r = 2'b01;
			14'b10001010101110: M1r = 2'b01;
			14'b11001010101110: M1r = 2'b01;
			14'b00011010101110: M1r = 2'b00;
			14'b01011010101110: M1r = 2'b00;
			14'b10011010101110: M1r = 2'b00;
			14'b11011010101110: M1r = 2'b01;
			14'b00101010101110: M1r = 2'b00;
			14'b01101010101110: M1r = 2'b00;
			14'b10101010101110: M1r = 2'b00;
			14'b11101010101110: M1r = 2'b00;
			14'b00111010101110: M1r = 2'b00;
			14'b01111010101110: M1r = 2'b00;
			14'b10111010101110: M1r = 2'b00;
			14'b11111010101110: M1r = 2'b00;
			14'b00001110101110: M1r = 2'b01;
			14'b01001110101110: M1r = 2'b01;
			14'b10001110101110: M1r = 2'b10;
			14'b11001110101110: M1r = 2'b10;
			14'b00011110101110: M1r = 2'b01;
			14'b01011110101110: M1r = 2'b01;
			14'b10011110101110: M1r = 2'b01;
			14'b11011110101110: M1r = 2'b01;
			14'b00101110101110: M1r = 2'b00;
			14'b01101110101110: M1r = 2'b01;
			14'b10101110101110: M1r = 2'b01;
			14'b11101110101110: M1r = 2'b01;
			14'b00111110101110: M1r = 2'b00;
			14'b01111110101110: M1r = 2'b00;
			14'b10111110101110: M1r = 2'b00;
			14'b11111110101110: M1r = 2'b00;
			14'b00000011101110: M1r = 2'b00;
			14'b01000011101110: M1r = 2'b00;
			14'b10000011101110: M1r = 2'b00;
			14'b11000011101110: M1r = 2'b00;
			14'b00010011101110: M1r = 2'b00;
			14'b01010011101110: M1r = 2'b00;
			14'b10010011101110: M1r = 2'b00;
			14'b11010011101110: M1r = 2'b00;
			14'b00100011101110: M1r = 2'b00;
			14'b01100011101110: M1r = 2'b00;
			14'b10100011101110: M1r = 2'b00;
			14'b11100011101110: M1r = 2'b00;
			14'b00110011101110: M1r = 2'b00;
			14'b01110011101110: M1r = 2'b00;
			14'b10110011101110: M1r = 2'b00;
			14'b11110011101110: M1r = 2'b00;
			14'b00000111101110: M1r = 2'b00;
			14'b01000111101110: M1r = 2'b00;
			14'b10000111101110: M1r = 2'b00;
			14'b11000111101110: M1r = 2'b00;
			14'b00010111101110: M1r = 2'b00;
			14'b01010111101110: M1r = 2'b00;
			14'b10010111101110: M1r = 2'b00;
			14'b11010111101110: M1r = 2'b00;
			14'b00100111101110: M1r = 2'b00;
			14'b01100111101110: M1r = 2'b00;
			14'b10100111101110: M1r = 2'b00;
			14'b11100111101110: M1r = 2'b00;
			14'b00110111101110: M1r = 2'b00;
			14'b01110111101110: M1r = 2'b00;
			14'b10110111101110: M1r = 2'b00;
			14'b11110111101110: M1r = 2'b00;
			14'b00001011101110: M1r = 2'b00;
			14'b01001011101110: M1r = 2'b00;
			14'b10001011101110: M1r = 2'b01;
			14'b11001011101110: M1r = 2'b01;
			14'b00011011101110: M1r = 2'b00;
			14'b01011011101110: M1r = 2'b00;
			14'b10011011101110: M1r = 2'b00;
			14'b11011011101110: M1r = 2'b00;
			14'b00101011101110: M1r = 2'b00;
			14'b01101011101110: M1r = 2'b00;
			14'b10101011101110: M1r = 2'b00;
			14'b11101011101110: M1r = 2'b00;
			14'b00111011101110: M1r = 2'b00;
			14'b01111011101110: M1r = 2'b00;
			14'b10111011101110: M1r = 2'b00;
			14'b11111011101110: M1r = 2'b00;
			14'b00001111101110: M1r = 2'b01;
			14'b01001111101110: M1r = 2'b01;
			14'b10001111101110: M1r = 2'b01;
			14'b11001111101110: M1r = 2'b01;
			14'b00011111101110: M1r = 2'b01;
			14'b01011111101110: M1r = 2'b01;
			14'b10011111101110: M1r = 2'b01;
			14'b11011111101110: M1r = 2'b01;
			14'b00101111101110: M1r = 2'b00;
			14'b01101111101110: M1r = 2'b00;
			14'b10101111101110: M1r = 2'b00;
			14'b11101111101110: M1r = 2'b01;
			14'b00111111101110: M1r = 2'b00;
			14'b01111111101110: M1r = 2'b00;
			14'b10111111101110: M1r = 2'b00;
			14'b11111111101110: M1r = 2'b00;
			14'b00000000111110: M1r = 2'b00;
			14'b01000000111110: M1r = 2'b00;
			14'b10000000111110: M1r = 2'b00;
			14'b11000000111110: M1r = 2'b01;
			14'b00010000111110: M1r = 2'b00;
			14'b01010000111110: M1r = 2'b00;
			14'b10010000111110: M1r = 2'b00;
			14'b11010000111110: M1r = 2'b00;
			14'b00100000111110: M1r = 2'b00;
			14'b01100000111110: M1r = 2'b00;
			14'b10100000111110: M1r = 2'b00;
			14'b11100000111110: M1r = 2'b00;
			14'b00110000111110: M1r = 2'b00;
			14'b01110000111110: M1r = 2'b00;
			14'b10110000111110: M1r = 2'b00;
			14'b11110000111110: M1r = 2'b00;
			14'b00000100111110: M1r = 2'b01;
			14'b01000100111110: M1r = 2'b01;
			14'b10000100111110: M1r = 2'b01;
			14'b11000100111110: M1r = 2'b01;
			14'b00010100111110: M1r = 2'b00;
			14'b01010100111110: M1r = 2'b00;
			14'b10010100111110: M1r = 2'b01;
			14'b11010100111110: M1r = 2'b01;
			14'b00100100111110: M1r = 2'b00;
			14'b01100100111110: M1r = 2'b00;
			14'b10100100111110: M1r = 2'b00;
			14'b11100100111110: M1r = 2'b00;
			14'b00110100111110: M1r = 2'b00;
			14'b01110100111110: M1r = 2'b00;
			14'b10110100111110: M1r = 2'b00;
			14'b11110100111110: M1r = 2'b00;
			14'b00001000111110: M1r = 2'b10;
			14'b01001000111110: M1r = 2'b10;
			14'b10001000111110: M1r = 2'b10;
			14'b11001000111110: M1r = 2'b10;
			14'b00011000111110: M1r = 2'b01;
			14'b01011000111110: M1r = 2'b01;
			14'b10011000111110: M1r = 2'b01;
			14'b11011000111110: M1r = 2'b10;
			14'b00101000111110: M1r = 2'b01;
			14'b01101000111110: M1r = 2'b01;
			14'b10101000111110: M1r = 2'b01;
			14'b11101000111110: M1r = 2'b01;
			14'b00111000111110: M1r = 2'b00;
			14'b01111000111110: M1r = 2'b00;
			14'b10111000111110: M1r = 2'b00;
			14'b11111000111110: M1r = 2'b01;
			14'b00001100111110: M1r = 2'b10;
			14'b01001100111110: M1r = 2'b10;
			14'b10001100111110: M1r = 2'b11;
			14'b11001100111110: M1r = 2'b11;
			14'b00011100111110: M1r = 2'b10;
			14'b01011100111110: M1r = 2'b10;
			14'b10011100111110: M1r = 2'b10;
			14'b11011100111110: M1r = 2'b10;
			14'b00101100111110: M1r = 2'b01;
			14'b01101100111110: M1r = 2'b01;
			14'b10101100111110: M1r = 2'b10;
			14'b11101100111110: M1r = 2'b10;
			14'b00111100111110: M1r = 2'b01;
			14'b01111100111110: M1r = 2'b01;
			14'b10111100111110: M1r = 2'b01;
			14'b11111100111110: M1r = 2'b01;
			14'b00000001111110: M1r = 2'b00;
			14'b01000001111110: M1r = 2'b00;
			14'b10000001111110: M1r = 2'b00;
			14'b11000001111110: M1r = 2'b00;
			14'b00010001111110: M1r = 2'b00;
			14'b01010001111110: M1r = 2'b00;
			14'b10010001111110: M1r = 2'b00;
			14'b11010001111110: M1r = 2'b00;
			14'b00100001111110: M1r = 2'b00;
			14'b01100001111110: M1r = 2'b00;
			14'b10100001111110: M1r = 2'b00;
			14'b11100001111110: M1r = 2'b00;
			14'b00110001111110: M1r = 2'b00;
			14'b01110001111110: M1r = 2'b00;
			14'b10110001111110: M1r = 2'b00;
			14'b11110001111110: M1r = 2'b00;
			14'b00000101111110: M1r = 2'b01;
			14'b01000101111110: M1r = 2'b01;
			14'b10000101111110: M1r = 2'b01;
			14'b11000101111110: M1r = 2'b01;
			14'b00010101111110: M1r = 2'b00;
			14'b01010101111110: M1r = 2'b00;
			14'b10010101111110: M1r = 2'b00;
			14'b11010101111110: M1r = 2'b01;
			14'b00100101111110: M1r = 2'b00;
			14'b01100101111110: M1r = 2'b00;
			14'b10100101111110: M1r = 2'b00;
			14'b11100101111110: M1r = 2'b00;
			14'b00110101111110: M1r = 2'b00;
			14'b01110101111110: M1r = 2'b00;
			14'b10110101111110: M1r = 2'b00;
			14'b11110101111110: M1r = 2'b00;
			14'b00001001111110: M1r = 2'b01;
			14'b01001001111110: M1r = 2'b01;
			14'b10001001111110: M1r = 2'b10;
			14'b11001001111110: M1r = 2'b10;
			14'b00011001111110: M1r = 2'b01;
			14'b01011001111110: M1r = 2'b01;
			14'b10011001111110: M1r = 2'b01;
			14'b11011001111110: M1r = 2'b01;
			14'b00101001111110: M1r = 2'b00;
			14'b01101001111110: M1r = 2'b00;
			14'b10101001111110: M1r = 2'b01;
			14'b11101001111110: M1r = 2'b01;
			14'b00111001111110: M1r = 2'b00;
			14'b01111001111110: M1r = 2'b00;
			14'b10111001111110: M1r = 2'b00;
			14'b11111001111110: M1r = 2'b00;
			14'b00001101111110: M1r = 2'b10;
			14'b01001101111110: M1r = 2'b10;
			14'b10001101111110: M1r = 2'b10;
			14'b11001101111110: M1r = 2'b10;
			14'b00011101111110: M1r = 2'b10;
			14'b01011101111110: M1r = 2'b10;
			14'b10011101111110: M1r = 2'b10;
			14'b11011101111110: M1r = 2'b10;
			14'b00101101111110: M1r = 2'b01;
			14'b01101101111110: M1r = 2'b01;
			14'b10101101111110: M1r = 2'b01;
			14'b11101101111110: M1r = 2'b10;
			14'b00111101111110: M1r = 2'b01;
			14'b01111101111110: M1r = 2'b01;
			14'b10111101111110: M1r = 2'b01;
			14'b11111101111110: M1r = 2'b01;
			14'b00000010111110: M1r = 2'b00;
			14'b01000010111110: M1r = 2'b00;
			14'b10000010111110: M1r = 2'b00;
			14'b11000010111110: M1r = 2'b00;
			14'b00010010111110: M1r = 2'b00;
			14'b01010010111110: M1r = 2'b00;
			14'b10010010111110: M1r = 2'b00;
			14'b11010010111110: M1r = 2'b00;
			14'b00100010111110: M1r = 2'b00;
			14'b01100010111110: M1r = 2'b00;
			14'b10100010111110: M1r = 2'b00;
			14'b11100010111110: M1r = 2'b00;
			14'b00110010111110: M1r = 2'b00;
			14'b01110010111110: M1r = 2'b00;
			14'b10110010111110: M1r = 2'b00;
			14'b11110010111110: M1r = 2'b00;
			14'b00000110111110: M1r = 2'b00;
			14'b01000110111110: M1r = 2'b00;
			14'b10000110111110: M1r = 2'b01;
			14'b11000110111110: M1r = 2'b01;
			14'b00010110111110: M1r = 2'b00;
			14'b01010110111110: M1r = 2'b00;
			14'b10010110111110: M1r = 2'b00;
			14'b11010110111110: M1r = 2'b00;
			14'b00100110111110: M1r = 2'b00;
			14'b01100110111110: M1r = 2'b00;
			14'b10100110111110: M1r = 2'b00;
			14'b11100110111110: M1r = 2'b00;
			14'b00110110111110: M1r = 2'b00;
			14'b01110110111110: M1r = 2'b00;
			14'b10110110111110: M1r = 2'b00;
			14'b11110110111110: M1r = 2'b00;
			14'b00001010111110: M1r = 2'b01;
			14'b01001010111110: M1r = 2'b01;
			14'b10001010111110: M1r = 2'b01;
			14'b11001010111110: M1r = 2'b01;
			14'b00011010111110: M1r = 2'b01;
			14'b01011010111110: M1r = 2'b01;
			14'b10011010111110: M1r = 2'b01;
			14'b11011010111110: M1r = 2'b01;
			14'b00101010111110: M1r = 2'b00;
			14'b01101010111110: M1r = 2'b00;
			14'b10101010111110: M1r = 2'b00;
			14'b11101010111110: M1r = 2'b01;
			14'b00111010111110: M1r = 2'b00;
			14'b01111010111110: M1r = 2'b00;
			14'b10111010111110: M1r = 2'b00;
			14'b11111010111110: M1r = 2'b00;
			14'b00001110111110: M1r = 2'b10;
			14'b01001110111110: M1r = 2'b10;
			14'b10001110111110: M1r = 2'b10;
			14'b11001110111110: M1r = 2'b10;
			14'b00011110111110: M1r = 2'b01;
			14'b01011110111110: M1r = 2'b01;
			14'b10011110111110: M1r = 2'b10;
			14'b11011110111110: M1r = 2'b10;
			14'b00101110111110: M1r = 2'b01;
			14'b01101110111110: M1r = 2'b01;
			14'b10101110111110: M1r = 2'b01;
			14'b11101110111110: M1r = 2'b01;
			14'b00111110111110: M1r = 2'b00;
			14'b01111110111110: M1r = 2'b00;
			14'b10111110111110: M1r = 2'b01;
			14'b11111110111110: M1r = 2'b01;
			14'b00000011111110: M1r = 2'b00;
			14'b01000011111110: M1r = 2'b00;
			14'b10000011111110: M1r = 2'b00;
			14'b11000011111110: M1r = 2'b00;
			14'b00010011111110: M1r = 2'b00;
			14'b01010011111110: M1r = 2'b00;
			14'b10010011111110: M1r = 2'b00;
			14'b11010011111110: M1r = 2'b00;
			14'b00100011111110: M1r = 2'b00;
			14'b01100011111110: M1r = 2'b00;
			14'b10100011111110: M1r = 2'b00;
			14'b11100011111110: M1r = 2'b00;
			14'b00110011111110: M1r = 2'b00;
			14'b01110011111110: M1r = 2'b00;
			14'b10110011111110: M1r = 2'b00;
			14'b11110011111110: M1r = 2'b00;
			14'b00000111111110: M1r = 2'b00;
			14'b01000111111110: M1r = 2'b00;
			14'b10000111111110: M1r = 2'b00;
			14'b11000111111110: M1r = 2'b00;
			14'b00010111111110: M1r = 2'b00;
			14'b01010111111110: M1r = 2'b00;
			14'b10010111111110: M1r = 2'b00;
			14'b11010111111110: M1r = 2'b00;
			14'b00100111111110: M1r = 2'b00;
			14'b01100111111110: M1r = 2'b00;
			14'b10100111111110: M1r = 2'b00;
			14'b11100111111110: M1r = 2'b00;
			14'b00110111111110: M1r = 2'b00;
			14'b01110111111110: M1r = 2'b00;
			14'b10110111111110: M1r = 2'b00;
			14'b11110111111110: M1r = 2'b00;
			14'b00001011111110: M1r = 2'b01;
			14'b01001011111110: M1r = 2'b01;
			14'b10001011111110: M1r = 2'b01;
			14'b11001011111110: M1r = 2'b01;
			14'b00011011111110: M1r = 2'b00;
			14'b01011011111110: M1r = 2'b00;
			14'b10011011111110: M1r = 2'b01;
			14'b11011011111110: M1r = 2'b01;
			14'b00101011111110: M1r = 2'b00;
			14'b01101011111110: M1r = 2'b00;
			14'b10101011111110: M1r = 2'b00;
			14'b11101011111110: M1r = 2'b00;
			14'b00111011111110: M1r = 2'b00;
			14'b01111011111110: M1r = 2'b00;
			14'b10111011111110: M1r = 2'b00;
			14'b11111011111110: M1r = 2'b00;
			14'b00001111111110: M1r = 2'b01;
			14'b01001111111110: M1r = 2'b10;
			14'b10001111111110: M1r = 2'b10;
			14'b11001111111110: M1r = 2'b10;
			14'b00011111111110: M1r = 2'b01;
			14'b01011111111110: M1r = 2'b01;
			14'b10011111111110: M1r = 2'b01;
			14'b11011111111110: M1r = 2'b01;
			14'b00101111111110: M1r = 2'b01;
			14'b01101111111110: M1r = 2'b01;
			14'b10101111111110: M1r = 2'b01;
			14'b11101111111110: M1r = 2'b01;
			14'b00111111111110: M1r = 2'b00;
			14'b01111111111110: M1r = 2'b00;
			14'b10111111111110: M1r = 2'b00;
			14'b11111111111110: M1r = 2'b01;
			14'b00000000000011: M1r = 2'b10;
			14'b01000000000011: M1r = 2'b10;
			14'b10000000000011: M1r = 2'b10;
			14'b11000000000011: M1r = 2'b11;
			14'b00010000000011: M1r = 2'b10;
			14'b01010000000011: M1r = 2'b10;
			14'b10010000000011: M1r = 2'b10;
			14'b11010000000011: M1r = 2'b10;
			14'b00100000000011: M1r = 2'b01;
			14'b01100000000011: M1r = 2'b01;
			14'b10100000000011: M1r = 2'b01;
			14'b11100000000011: M1r = 2'b10;
			14'b00110000000011: M1r = 2'b01;
			14'b01110000000011: M1r = 2'b01;
			14'b10110000000011: M1r = 2'b01;
			14'b11110000000011: M1r = 2'b01;
			14'b00000100000011: M1r = 2'b11;
			14'b01000100000011: M1r = 2'b11;
			14'b10000100000011: M1r = 2'b11;
			14'b11000100000011: M1r = 2'b11;
			14'b00010100000011: M1r = 2'b10;
			14'b01010100000011: M1r = 2'b10;
			14'b10010100000011: M1r = 2'b11;
			14'b11010100000011: M1r = 2'b11;
			14'b00100100000011: M1r = 2'b10;
			14'b01100100000011: M1r = 2'b10;
			14'b10100100000011: M1r = 2'b10;
			14'b11100100000011: M1r = 2'b10;
			14'b00110100000011: M1r = 2'b01;
			14'b01110100000011: M1r = 2'b10;
			14'b10110100000011: M1r = 2'b10;
			14'b11110100000011: M1r = 2'b10;
			14'b00001000000011: M1r = 2'b11;
			14'b01001000000011: M1r = 2'b11;
			14'b10001000000011: M1r = 2'b11;
			14'b11001000000011: M1r = 2'b11;
			14'b00011000000011: M1r = 2'b11;
			14'b01011000000011: M1r = 2'b11;
			14'b10011000000011: M1r = 2'b11;
			14'b11011000000011: M1r = 2'b11;
			14'b00101000000011: M1r = 2'b11;
			14'b01101000000011: M1r = 2'b11;
			14'b10101000000011: M1r = 2'b11;
			14'b11101000000011: M1r = 2'b11;
			14'b00111000000011: M1r = 2'b10;
			14'b01111000000011: M1r = 2'b10;
			14'b10111000000011: M1r = 2'b10;
			14'b11111000000011: M1r = 2'b11;
			14'b00001100000011: M1r = 2'b11;
			14'b01001100000011: M1r = 2'b11;
			14'b10001100000011: M1r = 2'b11;
			14'b11001100000011: M1r = 2'b11;
			14'b00011100000011: M1r = 2'b11;
			14'b01011100000011: M1r = 2'b11;
			14'b10011100000011: M1r = 2'b11;
			14'b11011100000011: M1r = 2'b11;
			14'b00101100000011: M1r = 2'b11;
			14'b01101100000011: M1r = 2'b11;
			14'b10101100000011: M1r = 2'b11;
			14'b11101100000011: M1r = 2'b11;
			14'b00111100000011: M1r = 2'b11;
			14'b01111100000011: M1r = 2'b11;
			14'b10111100000011: M1r = 2'b11;
			14'b11111100000011: M1r = 2'b11;
			14'b00000001000011: M1r = 2'b10;
			14'b01000001000011: M1r = 2'b10;
			14'b10000001000011: M1r = 2'b10;
			14'b11000001000011: M1r = 2'b10;
			14'b00010001000011: M1r = 2'b01;
			14'b01010001000011: M1r = 2'b01;
			14'b10010001000011: M1r = 2'b10;
			14'b11010001000011: M1r = 2'b10;
			14'b00100001000011: M1r = 2'b01;
			14'b01100001000011: M1r = 2'b01;
			14'b10100001000011: M1r = 2'b01;
			14'b11100001000011: M1r = 2'b01;
			14'b00110001000011: M1r = 2'b00;
			14'b01110001000011: M1r = 2'b01;
			14'b10110001000011: M1r = 2'b01;
			14'b11110001000011: M1r = 2'b01;
			14'b00000101000011: M1r = 2'b11;
			14'b01000101000011: M1r = 2'b11;
			14'b10000101000011: M1r = 2'b11;
			14'b11000101000011: M1r = 2'b11;
			14'b00010101000011: M1r = 2'b10;
			14'b01010101000011: M1r = 2'b10;
			14'b10010101000011: M1r = 2'b10;
			14'b11010101000011: M1r = 2'b11;
			14'b00100101000011: M1r = 2'b10;
			14'b01100101000011: M1r = 2'b10;
			14'b10100101000011: M1r = 2'b10;
			14'b11100101000011: M1r = 2'b10;
			14'b00110101000011: M1r = 2'b01;
			14'b01110101000011: M1r = 2'b01;
			14'b10110101000011: M1r = 2'b01;
			14'b11110101000011: M1r = 2'b10;
			14'b00001001000011: M1r = 2'b11;
			14'b01001001000011: M1r = 2'b11;
			14'b10001001000011: M1r = 2'b11;
			14'b11001001000011: M1r = 2'b11;
			14'b00011001000011: M1r = 2'b11;
			14'b01011001000011: M1r = 2'b11;
			14'b10011001000011: M1r = 2'b11;
			14'b11011001000011: M1r = 2'b11;
			14'b00101001000011: M1r = 2'b10;
			14'b01101001000011: M1r = 2'b10;
			14'b10101001000011: M1r = 2'b11;
			14'b11101001000011: M1r = 2'b11;
			14'b00111001000011: M1r = 2'b10;
			14'b01111001000011: M1r = 2'b10;
			14'b10111001000011: M1r = 2'b10;
			14'b11111001000011: M1r = 2'b10;
			14'b00001101000011: M1r = 2'b11;
			14'b01001101000011: M1r = 2'b11;
			14'b10001101000011: M1r = 2'b11;
			14'b11001101000011: M1r = 2'b11;
			14'b00011101000011: M1r = 2'b11;
			14'b01011101000011: M1r = 2'b11;
			14'b10011101000011: M1r = 2'b11;
			14'b11011101000011: M1r = 2'b11;
			14'b00101101000011: M1r = 2'b11;
			14'b01101101000011: M1r = 2'b11;
			14'b10101101000011: M1r = 2'b11;
			14'b11101101000011: M1r = 2'b11;
			14'b00111101000011: M1r = 2'b11;
			14'b01111101000011: M1r = 2'b11;
			14'b10111101000011: M1r = 2'b11;
			14'b11111101000011: M1r = 2'b11;
			14'b00000010000011: M1r = 2'b01;
			14'b01000010000011: M1r = 2'b10;
			14'b10000010000011: M1r = 2'b10;
			14'b11000010000011: M1r = 2'b10;
			14'b00010010000011: M1r = 2'b01;
			14'b01010010000011: M1r = 2'b01;
			14'b10010010000011: M1r = 2'b01;
			14'b11010010000011: M1r = 2'b01;
			14'b00100010000011: M1r = 2'b01;
			14'b01100010000011: M1r = 2'b01;
			14'b10100010000011: M1r = 2'b01;
			14'b11100010000011: M1r = 2'b01;
			14'b00110010000011: M1r = 2'b00;
			14'b01110010000011: M1r = 2'b00;
			14'b10110010000011: M1r = 2'b00;
			14'b11110010000011: M1r = 2'b01;
			14'b00000110000011: M1r = 2'b10;
			14'b01000110000011: M1r = 2'b10;
			14'b10000110000011: M1r = 2'b11;
			14'b11000110000011: M1r = 2'b11;
			14'b00010110000011: M1r = 2'b10;
			14'b01010110000011: M1r = 2'b10;
			14'b10010110000011: M1r = 2'b10;
			14'b11010110000011: M1r = 2'b10;
			14'b00100110000011: M1r = 2'b01;
			14'b01100110000011: M1r = 2'b01;
			14'b10100110000011: M1r = 2'b10;
			14'b11100110000011: M1r = 2'b10;
			14'b00110110000011: M1r = 2'b01;
			14'b01110110000011: M1r = 2'b01;
			14'b10110110000011: M1r = 2'b01;
			14'b11110110000011: M1r = 2'b01;
			14'b00001010000011: M1r = 2'b11;
			14'b01001010000011: M1r = 2'b11;
			14'b10001010000011: M1r = 2'b11;
			14'b11001010000011: M1r = 2'b11;
			14'b00011010000011: M1r = 2'b11;
			14'b01011010000011: M1r = 2'b11;
			14'b10011010000011: M1r = 2'b11;
			14'b11011010000011: M1r = 2'b11;
			14'b00101010000011: M1r = 2'b10;
			14'b01101010000011: M1r = 2'b10;
			14'b10101010000011: M1r = 2'b10;
			14'b11101010000011: M1r = 2'b11;
			14'b00111010000011: M1r = 2'b10;
			14'b01111010000011: M1r = 2'b10;
			14'b10111010000011: M1r = 2'b10;
			14'b11111010000011: M1r = 2'b10;
			14'b00001110000011: M1r = 2'b11;
			14'b01001110000011: M1r = 2'b11;
			14'b10001110000011: M1r = 2'b11;
			14'b11001110000011: M1r = 2'b11;
			14'b00011110000011: M1r = 2'b11;
			14'b01011110000011: M1r = 2'b11;
			14'b10011110000011: M1r = 2'b11;
			14'b11011110000011: M1r = 2'b11;
			14'b00101110000011: M1r = 2'b11;
			14'b01101110000011: M1r = 2'b11;
			14'b10101110000011: M1r = 2'b11;
			14'b11101110000011: M1r = 2'b11;
			14'b00111110000011: M1r = 2'b10;
			14'b01111110000011: M1r = 2'b10;
			14'b10111110000011: M1r = 2'b11;
			14'b11111110000011: M1r = 2'b11;
			14'b00000011000011: M1r = 2'b01;
			14'b01000011000011: M1r = 2'b01;
			14'b10000011000011: M1r = 2'b10;
			14'b11000011000011: M1r = 2'b10;
			14'b00010011000011: M1r = 2'b01;
			14'b01010011000011: M1r = 2'b01;
			14'b10010011000011: M1r = 2'b01;
			14'b11010011000011: M1r = 2'b01;
			14'b00100011000011: M1r = 2'b00;
			14'b01100011000011: M1r = 2'b00;
			14'b10100011000011: M1r = 2'b01;
			14'b11100011000011: M1r = 2'b01;
			14'b00110011000011: M1r = 2'b00;
			14'b01110011000011: M1r = 2'b00;
			14'b10110011000011: M1r = 2'b00;
			14'b11110011000011: M1r = 2'b00;
			14'b00000111000011: M1r = 2'b10;
			14'b01000111000011: M1r = 2'b10;
			14'b10000111000011: M1r = 2'b10;
			14'b11000111000011: M1r = 2'b10;
			14'b00010111000011: M1r = 2'b01;
			14'b01010111000011: M1r = 2'b10;
			14'b10010111000011: M1r = 2'b10;
			14'b11010111000011: M1r = 2'b10;
			14'b00100111000011: M1r = 2'b01;
			14'b01100111000011: M1r = 2'b01;
			14'b10100111000011: M1r = 2'b01;
			14'b11100111000011: M1r = 2'b01;
			14'b00110111000011: M1r = 2'b01;
			14'b01110111000011: M1r = 2'b01;
			14'b10110111000011: M1r = 2'b01;
			14'b11110111000011: M1r = 2'b01;
			14'b00001011000011: M1r = 2'b11;
			14'b01001011000011: M1r = 2'b11;
			14'b10001011000011: M1r = 2'b11;
			14'b11001011000011: M1r = 2'b11;
			14'b00011011000011: M1r = 2'b10;
			14'b01011011000011: M1r = 2'b10;
			14'b10011011000011: M1r = 2'b11;
			14'b11011011000011: M1r = 2'b11;
			14'b00101011000011: M1r = 2'b10;
			14'b01101011000011: M1r = 2'b10;
			14'b10101011000011: M1r = 2'b10;
			14'b11101011000011: M1r = 2'b10;
			14'b00111011000011: M1r = 2'b01;
			14'b01111011000011: M1r = 2'b01;
			14'b10111011000011: M1r = 2'b10;
			14'b11111011000011: M1r = 2'b10;
			14'b00001111000011: M1r = 2'b11;
			14'b01001111000011: M1r = 2'b11;
			14'b10001111000011: M1r = 2'b11;
			14'b11001111000011: M1r = 2'b11;
			14'b00011111000011: M1r = 2'b11;
			14'b01011111000011: M1r = 2'b11;
			14'b10011111000011: M1r = 2'b11;
			14'b11011111000011: M1r = 2'b11;
			14'b00101111000011: M1r = 2'b11;
			14'b01101111000011: M1r = 2'b11;
			14'b10101111000011: M1r = 2'b11;
			14'b11101111000011: M1r = 2'b11;
			14'b00111111000011: M1r = 2'b10;
			14'b01111111000011: M1r = 2'b10;
			14'b10111111000011: M1r = 2'b10;
			14'b11111111000011: M1r = 2'b11;
			14'b00000000010011: M1r = 2'b10;
			14'b01000000010011: M1r = 2'b11;
			14'b10000000010011: M1r = 2'b11;
			14'b11000000010011: M1r = 2'b11;
			14'b00010000010011: M1r = 2'b10;
			14'b01010000010011: M1r = 2'b10;
			14'b10010000010011: M1r = 2'b10;
			14'b11010000010011: M1r = 2'b10;
			14'b00100000010011: M1r = 2'b10;
			14'b01100000010011: M1r = 2'b10;
			14'b10100000010011: M1r = 2'b10;
			14'b11100000010011: M1r = 2'b10;
			14'b00110000010011: M1r = 2'b01;
			14'b01110000010011: M1r = 2'b01;
			14'b10110000010011: M1r = 2'b01;
			14'b11110000010011: M1r = 2'b10;
			14'b00000100010011: M1r = 2'b11;
			14'b01000100010011: M1r = 2'b11;
			14'b10000100010011: M1r = 2'b11;
			14'b11000100010011: M1r = 2'b11;
			14'b00010100010011: M1r = 2'b11;
			14'b01010100010011: M1r = 2'b11;
			14'b10010100010011: M1r = 2'b11;
			14'b11010100010011: M1r = 2'b11;
			14'b00100100010011: M1r = 2'b10;
			14'b01100100010011: M1r = 2'b10;
			14'b10100100010011: M1r = 2'b11;
			14'b11100100010011: M1r = 2'b11;
			14'b00110100010011: M1r = 2'b10;
			14'b01110100010011: M1r = 2'b10;
			14'b10110100010011: M1r = 2'b10;
			14'b11110100010011: M1r = 2'b10;
			14'b00001000010011: M1r = 2'b11;
			14'b01001000010011: M1r = 2'b11;
			14'b10001000010011: M1r = 2'b11;
			14'b11001000010011: M1r = 2'b11;
			14'b00011000010011: M1r = 2'b11;
			14'b01011000010011: M1r = 2'b11;
			14'b10011000010011: M1r = 2'b11;
			14'b11011000010011: M1r = 2'b11;
			14'b00101000010011: M1r = 2'b11;
			14'b01101000010011: M1r = 2'b11;
			14'b10101000010011: M1r = 2'b11;
			14'b11101000010011: M1r = 2'b11;
			14'b00111000010011: M1r = 2'b11;
			14'b01111000010011: M1r = 2'b11;
			14'b10111000010011: M1r = 2'b11;
			14'b11111000010011: M1r = 2'b11;
			14'b00001100010011: M1r = 2'b11;
			14'b01001100010011: M1r = 2'b11;
			14'b10001100010011: M1r = 2'b11;
			14'b11001100010011: M1r = 2'b11;
			14'b00011100010011: M1r = 2'b11;
			14'b01011100010011: M1r = 2'b11;
			14'b10011100010011: M1r = 2'b11;
			14'b11011100010011: M1r = 2'b11;
			14'b00101100010011: M1r = 2'b11;
			14'b01101100010011: M1r = 2'b11;
			14'b10101100010011: M1r = 2'b11;
			14'b11101100010011: M1r = 2'b11;
			14'b00111100010011: M1r = 2'b11;
			14'b01111100010011: M1r = 2'b11;
			14'b10111100010011: M1r = 2'b11;
			14'b11111100010011: M1r = 2'b11;
			14'b00000001010011: M1r = 2'b10;
			14'b01000001010011: M1r = 2'b10;
			14'b10000001010011: M1r = 2'b11;
			14'b11000001010011: M1r = 2'b11;
			14'b00010001010011: M1r = 2'b10;
			14'b01010001010011: M1r = 2'b10;
			14'b10010001010011: M1r = 2'b10;
			14'b11010001010011: M1r = 2'b10;
			14'b00100001010011: M1r = 2'b01;
			14'b01100001010011: M1r = 2'b01;
			14'b10100001010011: M1r = 2'b10;
			14'b11100001010011: M1r = 2'b10;
			14'b00110001010011: M1r = 2'b01;
			14'b01110001010011: M1r = 2'b01;
			14'b10110001010011: M1r = 2'b01;
			14'b11110001010011: M1r = 2'b01;
			14'b00000101010011: M1r = 2'b11;
			14'b01000101010011: M1r = 2'b11;
			14'b10000101010011: M1r = 2'b11;
			14'b11000101010011: M1r = 2'b11;
			14'b00010101010011: M1r = 2'b10;
			14'b01010101010011: M1r = 2'b11;
			14'b10010101010011: M1r = 2'b11;
			14'b11010101010011: M1r = 2'b11;
			14'b00100101010011: M1r = 2'b10;
			14'b01100101010011: M1r = 2'b10;
			14'b10100101010011: M1r = 2'b10;
			14'b11100101010011: M1r = 2'b10;
			14'b00110101010011: M1r = 2'b10;
			14'b01110101010011: M1r = 2'b10;
			14'b10110101010011: M1r = 2'b10;
			14'b11110101010011: M1r = 2'b10;
			14'b00001001010011: M1r = 2'b11;
			14'b01001001010011: M1r = 2'b11;
			14'b10001001010011: M1r = 2'b11;
			14'b11001001010011: M1r = 2'b11;
			14'b00011001010011: M1r = 2'b11;
			14'b01011001010011: M1r = 2'b11;
			14'b10011001010011: M1r = 2'b11;
			14'b11011001010011: M1r = 2'b11;
			14'b00101001010011: M1r = 2'b11;
			14'b01101001010011: M1r = 2'b11;
			14'b10101001010011: M1r = 2'b11;
			14'b11101001010011: M1r = 2'b11;
			14'b00111001010011: M1r = 2'b10;
			14'b01111001010011: M1r = 2'b10;
			14'b10111001010011: M1r = 2'b11;
			14'b11111001010011: M1r = 2'b11;
			14'b00001101010011: M1r = 2'b11;
			14'b01001101010011: M1r = 2'b11;
			14'b10001101010011: M1r = 2'b11;
			14'b11001101010011: M1r = 2'b11;
			14'b00011101010011: M1r = 2'b11;
			14'b01011101010011: M1r = 2'b11;
			14'b10011101010011: M1r = 2'b11;
			14'b11011101010011: M1r = 2'b11;
			14'b00101101010011: M1r = 2'b11;
			14'b01101101010011: M1r = 2'b11;
			14'b10101101010011: M1r = 2'b11;
			14'b11101101010011: M1r = 2'b11;
			14'b00111101010011: M1r = 2'b11;
			14'b01111101010011: M1r = 2'b11;
			14'b10111101010011: M1r = 2'b11;
			14'b11111101010011: M1r = 2'b11;
			14'b00000010010011: M1r = 2'b10;
			14'b01000010010011: M1r = 2'b10;
			14'b10000010010011: M1r = 2'b10;
			14'b11000010010011: M1r = 2'b10;
			14'b00010010010011: M1r = 2'b01;
			14'b01010010010011: M1r = 2'b10;
			14'b10010010010011: M1r = 2'b10;
			14'b11010010010011: M1r = 2'b10;
			14'b00100010010011: M1r = 2'b01;
			14'b01100010010011: M1r = 2'b01;
			14'b10100010010011: M1r = 2'b01;
			14'b11100010010011: M1r = 2'b01;
			14'b00110010010011: M1r = 2'b01;
			14'b01110010010011: M1r = 2'b01;
			14'b10110010010011: M1r = 2'b01;
			14'b11110010010011: M1r = 2'b01;
			14'b00000110010011: M1r = 2'b11;
			14'b01000110010011: M1r = 2'b11;
			14'b10000110010011: M1r = 2'b11;
			14'b11000110010011: M1r = 2'b11;
			14'b00010110010011: M1r = 2'b10;
			14'b01010110010011: M1r = 2'b10;
			14'b10010110010011: M1r = 2'b11;
			14'b11010110010011: M1r = 2'b11;
			14'b00100110010011: M1r = 2'b10;
			14'b01100110010011: M1r = 2'b10;
			14'b10100110010011: M1r = 2'b10;
			14'b11100110010011: M1r = 2'b10;
			14'b00110110010011: M1r = 2'b01;
			14'b01110110010011: M1r = 2'b01;
			14'b10110110010011: M1r = 2'b10;
			14'b11110110010011: M1r = 2'b10;
			14'b00001010010011: M1r = 2'b11;
			14'b01001010010011: M1r = 2'b11;
			14'b10001010010011: M1r = 2'b11;
			14'b11001010010011: M1r = 2'b11;
			14'b00011010010011: M1r = 2'b11;
			14'b01011010010011: M1r = 2'b11;
			14'b10011010010011: M1r = 2'b11;
			14'b11011010010011: M1r = 2'b11;
			14'b00101010010011: M1r = 2'b10;
			14'b01101010010011: M1r = 2'b11;
			14'b10101010010011: M1r = 2'b11;
			14'b11101010010011: M1r = 2'b11;
			14'b00111010010011: M1r = 2'b10;
			14'b01111010010011: M1r = 2'b10;
			14'b10111010010011: M1r = 2'b10;
			14'b11111010010011: M1r = 2'b10;
			14'b00001110010011: M1r = 2'b11;
			14'b01001110010011: M1r = 2'b11;
			14'b10001110010011: M1r = 2'b11;
			14'b11001110010011: M1r = 2'b11;
			14'b00011110010011: M1r = 2'b11;
			14'b01011110010011: M1r = 2'b11;
			14'b10011110010011: M1r = 2'b11;
			14'b11011110010011: M1r = 2'b11;
			14'b00101110010011: M1r = 2'b11;
			14'b01101110010011: M1r = 2'b11;
			14'b10101110010011: M1r = 2'b11;
			14'b11101110010011: M1r = 2'b11;
			14'b00111110010011: M1r = 2'b11;
			14'b01111110010011: M1r = 2'b11;
			14'b10111110010011: M1r = 2'b11;
			14'b11111110010011: M1r = 2'b11;
			14'b00000011010011: M1r = 2'b10;
			14'b01000011010011: M1r = 2'b10;
			14'b10000011010011: M1r = 2'b10;
			14'b11000011010011: M1r = 2'b10;
			14'b00010011010011: M1r = 2'b01;
			14'b01010011010011: M1r = 2'b01;
			14'b10010011010011: M1r = 2'b01;
			14'b11010011010011: M1r = 2'b10;
			14'b00100011010011: M1r = 2'b01;
			14'b01100011010011: M1r = 2'b01;
			14'b10100011010011: M1r = 2'b01;
			14'b11100011010011: M1r = 2'b01;
			14'b00110011010011: M1r = 2'b00;
			14'b01110011010011: M1r = 2'b00;
			14'b10110011010011: M1r = 2'b01;
			14'b11110011010011: M1r = 2'b01;
			14'b00000111010011: M1r = 2'b10;
			14'b01000111010011: M1r = 2'b11;
			14'b10000111010011: M1r = 2'b11;
			14'b11000111010011: M1r = 2'b11;
			14'b00010111010011: M1r = 2'b10;
			14'b01010111010011: M1r = 2'b10;
			14'b10010111010011: M1r = 2'b10;
			14'b11010111010011: M1r = 2'b10;
			14'b00100111010011: M1r = 2'b01;
			14'b01100111010011: M1r = 2'b10;
			14'b10100111010011: M1r = 2'b10;
			14'b11100111010011: M1r = 2'b10;
			14'b00110111010011: M1r = 2'b01;
			14'b01110111010011: M1r = 2'b01;
			14'b10110111010011: M1r = 2'b01;
			14'b11110111010011: M1r = 2'b01;
			14'b00001011010011: M1r = 2'b11;
			14'b01001011010011: M1r = 2'b11;
			14'b10001011010011: M1r = 2'b11;
			14'b11001011010011: M1r = 2'b11;
			14'b00011011010011: M1r = 2'b11;
			14'b01011011010011: M1r = 2'b11;
			14'b10011011010011: M1r = 2'b11;
			14'b11011011010011: M1r = 2'b11;
			14'b00101011010011: M1r = 2'b10;
			14'b01101011010011: M1r = 2'b10;
			14'b10101011010011: M1r = 2'b11;
			14'b11101011010011: M1r = 2'b11;
			14'b00111011010011: M1r = 2'b10;
			14'b01111011010011: M1r = 2'b10;
			14'b10111011010011: M1r = 2'b10;
			14'b11111011010011: M1r = 2'b10;
			14'b00001111010011: M1r = 2'b11;
			14'b01001111010011: M1r = 2'b11;
			14'b10001111010011: M1r = 2'b11;
			14'b11001111010011: M1r = 2'b11;
			14'b00011111010011: M1r = 2'b11;
			14'b01011111010011: M1r = 2'b11;
			14'b10011111010011: M1r = 2'b11;
			14'b11011111010011: M1r = 2'b11;
			14'b00101111010011: M1r = 2'b11;
			14'b01101111010011: M1r = 2'b11;
			14'b10101111010011: M1r = 2'b11;
			14'b11101111010011: M1r = 2'b11;
			14'b00111111010011: M1r = 2'b10;
			14'b01111111010011: M1r = 2'b11;
			14'b10111111010011: M1r = 2'b11;
			14'b11111111010011: M1r = 2'b11;
			14'b00000000100011: M1r = 2'b11;
			14'b01000000100011: M1r = 2'b11;
			14'b10000000100011: M1r = 2'b11;
			14'b11000000100011: M1r = 2'b11;
			14'b00010000100011: M1r = 2'b10;
			14'b01010000100011: M1r = 2'b11;
			14'b10010000100011: M1r = 2'b11;
			14'b11010000100011: M1r = 2'b11;
			14'b00100000100011: M1r = 2'b10;
			14'b01100000100011: M1r = 2'b10;
			14'b10100000100011: M1r = 2'b10;
			14'b11100000100011: M1r = 2'b10;
			14'b00110000100011: M1r = 2'b01;
			14'b01110000100011: M1r = 2'b10;
			14'b10110000100011: M1r = 2'b10;
			14'b11110000100011: M1r = 2'b10;
			14'b00000100100011: M1r = 2'b11;
			14'b01000100100011: M1r = 2'b11;
			14'b10000100100011: M1r = 2'b11;
			14'b11000100100011: M1r = 2'b11;
			14'b00010100100011: M1r = 2'b11;
			14'b01010100100011: M1r = 2'b11;
			14'b10010100100011: M1r = 2'b11;
			14'b11010100100011: M1r = 2'b11;
			14'b00100100100011: M1r = 2'b11;
			14'b01100100100011: M1r = 2'b11;
			14'b10100100100011: M1r = 2'b11;
			14'b11100100100011: M1r = 2'b11;
			14'b00110100100011: M1r = 2'b10;
			14'b01110100100011: M1r = 2'b10;
			14'b10110100100011: M1r = 2'b11;
			14'b11110100100011: M1r = 2'b11;
			14'b00001000100011: M1r = 2'b11;
			14'b01001000100011: M1r = 2'b11;
			14'b10001000100011: M1r = 2'b11;
			14'b11001000100011: M1r = 2'b11;
			14'b00011000100011: M1r = 2'b11;
			14'b01011000100011: M1r = 2'b11;
			14'b10011000100011: M1r = 2'b11;
			14'b11011000100011: M1r = 2'b11;
			14'b00101000100011: M1r = 2'b11;
			14'b01101000100011: M1r = 2'b11;
			14'b10101000100011: M1r = 2'b11;
			14'b11101000100011: M1r = 2'b11;
			14'b00111000100011: M1r = 2'b11;
			14'b01111000100011: M1r = 2'b11;
			14'b10111000100011: M1r = 2'b11;
			14'b11111000100011: M1r = 2'b11;
			14'b00001100100011: M1r = 2'b11;
			14'b01001100100011: M1r = 2'b11;
			14'b10001100100011: M1r = 2'b11;
			14'b11001100100011: M1r = 2'b11;
			14'b00011100100011: M1r = 2'b11;
			14'b01011100100011: M1r = 2'b11;
			14'b10011100100011: M1r = 2'b11;
			14'b11011100100011: M1r = 2'b11;
			14'b00101100100011: M1r = 2'b11;
			14'b01101100100011: M1r = 2'b11;
			14'b10101100100011: M1r = 2'b11;
			14'b11101100100011: M1r = 2'b11;
			14'b00111100100011: M1r = 2'b11;
			14'b01111100100011: M1r = 2'b11;
			14'b10111100100011: M1r = 2'b11;
			14'b11111100100011: M1r = 2'b11;
			14'b00000001100011: M1r = 2'b11;
			14'b01000001100011: M1r = 2'b11;
			14'b10000001100011: M1r = 2'b11;
			14'b11000001100011: M1r = 2'b11;
			14'b00010001100011: M1r = 2'b10;
			14'b01010001100011: M1r = 2'b10;
			14'b10010001100011: M1r = 2'b10;
			14'b11010001100011: M1r = 2'b11;
			14'b00100001100011: M1r = 2'b10;
			14'b01100001100011: M1r = 2'b10;
			14'b10100001100011: M1r = 2'b10;
			14'b11100001100011: M1r = 2'b10;
			14'b00110001100011: M1r = 2'b01;
			14'b01110001100011: M1r = 2'b01;
			14'b10110001100011: M1r = 2'b10;
			14'b11110001100011: M1r = 2'b10;
			14'b00000101100011: M1r = 2'b11;
			14'b01000101100011: M1r = 2'b11;
			14'b10000101100011: M1r = 2'b11;
			14'b11000101100011: M1r = 2'b11;
			14'b00010101100011: M1r = 2'b11;
			14'b01010101100011: M1r = 2'b11;
			14'b10010101100011: M1r = 2'b11;
			14'b11010101100011: M1r = 2'b11;
			14'b00100101100011: M1r = 2'b10;
			14'b01100101100011: M1r = 2'b11;
			14'b10100101100011: M1r = 2'b11;
			14'b11100101100011: M1r = 2'b11;
			14'b00110101100011: M1r = 2'b10;
			14'b01110101100011: M1r = 2'b10;
			14'b10110101100011: M1r = 2'b10;
			14'b11110101100011: M1r = 2'b10;
			14'b00001001100011: M1r = 2'b11;
			14'b01001001100011: M1r = 2'b11;
			14'b10001001100011: M1r = 2'b11;
			14'b11001001100011: M1r = 2'b11;
			14'b00011001100011: M1r = 2'b11;
			14'b01011001100011: M1r = 2'b11;
			14'b10011001100011: M1r = 2'b11;
			14'b11011001100011: M1r = 2'b11;
			14'b00101001100011: M1r = 2'b11;
			14'b01101001100011: M1r = 2'b11;
			14'b10101001100011: M1r = 2'b11;
			14'b11101001100011: M1r = 2'b11;
			14'b00111001100011: M1r = 2'b11;
			14'b01111001100011: M1r = 2'b11;
			14'b10111001100011: M1r = 2'b11;
			14'b11111001100011: M1r = 2'b11;
			14'b00001101100011: M1r = 2'b11;
			14'b01001101100011: M1r = 2'b11;
			14'b10001101100011: M1r = 2'b11;
			14'b11001101100011: M1r = 2'b11;
			14'b00011101100011: M1r = 2'b11;
			14'b01011101100011: M1r = 2'b11;
			14'b10011101100011: M1r = 2'b11;
			14'b11011101100011: M1r = 2'b11;
			14'b00101101100011: M1r = 2'b11;
			14'b01101101100011: M1r = 2'b11;
			14'b10101101100011: M1r = 2'b11;
			14'b11101101100011: M1r = 2'b11;
			14'b00111101100011: M1r = 2'b11;
			14'b01111101100011: M1r = 2'b11;
			14'b10111101100011: M1r = 2'b11;
			14'b11111101100011: M1r = 2'b11;
			14'b00000010100011: M1r = 2'b10;
			14'b01000010100011: M1r = 2'b11;
			14'b10000010100011: M1r = 2'b11;
			14'b11000010100011: M1r = 2'b11;
			14'b00010010100011: M1r = 2'b10;
			14'b01010010100011: M1r = 2'b10;
			14'b10010010100011: M1r = 2'b10;
			14'b11010010100011: M1r = 2'b10;
			14'b00100010100011: M1r = 2'b01;
			14'b01100010100011: M1r = 2'b10;
			14'b10100010100011: M1r = 2'b10;
			14'b11100010100011: M1r = 2'b10;
			14'b00110010100011: M1r = 2'b01;
			14'b01110010100011: M1r = 2'b01;
			14'b10110010100011: M1r = 2'b01;
			14'b11110010100011: M1r = 2'b01;
			14'b00000110100011: M1r = 2'b11;
			14'b01000110100011: M1r = 2'b11;
			14'b10000110100011: M1r = 2'b11;
			14'b11000110100011: M1r = 2'b11;
			14'b00010110100011: M1r = 2'b11;
			14'b01010110100011: M1r = 2'b11;
			14'b10010110100011: M1r = 2'b11;
			14'b11010110100011: M1r = 2'b11;
			14'b00100110100011: M1r = 2'b10;
			14'b01100110100011: M1r = 2'b10;
			14'b10100110100011: M1r = 2'b10;
			14'b11100110100011: M1r = 2'b11;
			14'b00110110100011: M1r = 2'b10;
			14'b01110110100011: M1r = 2'b10;
			14'b10110110100011: M1r = 2'b10;
			14'b11110110100011: M1r = 2'b10;
			14'b00001010100011: M1r = 2'b11;
			14'b01001010100011: M1r = 2'b11;
			14'b10001010100011: M1r = 2'b11;
			14'b11001010100011: M1r = 2'b11;
			14'b00011010100011: M1r = 2'b11;
			14'b01011010100011: M1r = 2'b11;
			14'b10011010100011: M1r = 2'b11;
			14'b11011010100011: M1r = 2'b11;
			14'b00101010100011: M1r = 2'b11;
			14'b01101010100011: M1r = 2'b11;
			14'b10101010100011: M1r = 2'b11;
			14'b11101010100011: M1r = 2'b11;
			14'b00111010100011: M1r = 2'b10;
			14'b01111010100011: M1r = 2'b11;
			14'b10111010100011: M1r = 2'b11;
			14'b11111010100011: M1r = 2'b11;
			14'b00001110100011: M1r = 2'b11;
			14'b01001110100011: M1r = 2'b11;
			14'b10001110100011: M1r = 2'b11;
			14'b11001110100011: M1r = 2'b11;
			14'b00011110100011: M1r = 2'b11;
			14'b01011110100011: M1r = 2'b11;
			14'b10011110100011: M1r = 2'b11;
			14'b11011110100011: M1r = 2'b11;
			14'b00101110100011: M1r = 2'b11;
			14'b01101110100011: M1r = 2'b11;
			14'b10101110100011: M1r = 2'b11;
			14'b11101110100011: M1r = 2'b11;
			14'b00111110100011: M1r = 2'b11;
			14'b01111110100011: M1r = 2'b11;
			14'b10111110100011: M1r = 2'b11;
			14'b11111110100011: M1r = 2'b11;
			14'b00000011100011: M1r = 2'b10;
			14'b01000011100011: M1r = 2'b10;
			14'b10000011100011: M1r = 2'b10;
			14'b11000011100011: M1r = 2'b11;
			14'b00010011100011: M1r = 2'b10;
			14'b01010011100011: M1r = 2'b10;
			14'b10010011100011: M1r = 2'b10;
			14'b11010011100011: M1r = 2'b10;
			14'b00100011100011: M1r = 2'b01;
			14'b01100011100011: M1r = 2'b01;
			14'b10100011100011: M1r = 2'b01;
			14'b11100011100011: M1r = 2'b10;
			14'b00110011100011: M1r = 2'b01;
			14'b01110011100011: M1r = 2'b01;
			14'b10110011100011: M1r = 2'b01;
			14'b11110011100011: M1r = 2'b01;
			14'b00000111100011: M1r = 2'b11;
			14'b01000111100011: M1r = 2'b11;
			14'b10000111100011: M1r = 2'b11;
			14'b11000111100011: M1r = 2'b11;
			14'b00010111100011: M1r = 2'b10;
			14'b01010111100011: M1r = 2'b11;
			14'b10010111100011: M1r = 2'b11;
			14'b11010111100011: M1r = 2'b11;
			14'b00100111100011: M1r = 2'b10;
			14'b01100111100011: M1r = 2'b10;
			14'b10100111100011: M1r = 2'b10;
			14'b11100111100011: M1r = 2'b10;
			14'b00110111100011: M1r = 2'b01;
			14'b01110111100011: M1r = 2'b10;
			14'b10110111100011: M1r = 2'b10;
			14'b11110111100011: M1r = 2'b10;
			14'b00001011100011: M1r = 2'b11;
			14'b01001011100011: M1r = 2'b11;
			14'b10001011100011: M1r = 2'b11;
			14'b11001011100011: M1r = 2'b11;
			14'b00011011100011: M1r = 2'b11;
			14'b01011011100011: M1r = 2'b11;
			14'b10011011100011: M1r = 2'b11;
			14'b11011011100011: M1r = 2'b11;
			14'b00101011100011: M1r = 2'b11;
			14'b01101011100011: M1r = 2'b11;
			14'b10101011100011: M1r = 2'b11;
			14'b11101011100011: M1r = 2'b11;
			14'b00111011100011: M1r = 2'b10;
			14'b01111011100011: M1r = 2'b10;
			14'b10111011100011: M1r = 2'b10;
			14'b11111011100011: M1r = 2'b11;
			14'b00001111100011: M1r = 2'b11;
			14'b01001111100011: M1r = 2'b11;
			14'b10001111100011: M1r = 2'b11;
			14'b11001111100011: M1r = 2'b11;
			14'b00011111100011: M1r = 2'b11;
			14'b01011111100011: M1r = 2'b11;
			14'b10011111100011: M1r = 2'b11;
			14'b11011111100011: M1r = 2'b11;
			14'b00101111100011: M1r = 2'b11;
			14'b01101111100011: M1r = 2'b11;
			14'b10101111100011: M1r = 2'b11;
			14'b11101111100011: M1r = 2'b11;
			14'b00111111100011: M1r = 2'b11;
			14'b01111111100011: M1r = 2'b11;
			14'b10111111100011: M1r = 2'b11;
			14'b11111111100011: M1r = 2'b11;
			14'b00000000110011: M1r = 2'b11;
			14'b01000000110011: M1r = 2'b11;
			14'b10000000110011: M1r = 2'b11;
			14'b11000000110011: M1r = 2'b11;
			14'b00010000110011: M1r = 2'b11;
			14'b01010000110011: M1r = 2'b11;
			14'b10010000110011: M1r = 2'b11;
			14'b11010000110011: M1r = 2'b11;
			14'b00100000110011: M1r = 2'b10;
			14'b01100000110011: M1r = 2'b11;
			14'b10100000110011: M1r = 2'b11;
			14'b11100000110011: M1r = 2'b11;
			14'b00110000110011: M1r = 2'b10;
			14'b01110000110011: M1r = 2'b10;
			14'b10110000110011: M1r = 2'b10;
			14'b11110000110011: M1r = 2'b10;
			14'b00000100110011: M1r = 2'b11;
			14'b01000100110011: M1r = 2'b11;
			14'b10000100110011: M1r = 2'b11;
			14'b11000100110011: M1r = 2'b11;
			14'b00010100110011: M1r = 2'b11;
			14'b01010100110011: M1r = 2'b11;
			14'b10010100110011: M1r = 2'b11;
			14'b11010100110011: M1r = 2'b11;
			14'b00100100110011: M1r = 2'b11;
			14'b01100100110011: M1r = 2'b11;
			14'b10100100110011: M1r = 2'b11;
			14'b11100100110011: M1r = 2'b11;
			14'b00110100110011: M1r = 2'b11;
			14'b01110100110011: M1r = 2'b11;
			14'b10110100110011: M1r = 2'b11;
			14'b11110100110011: M1r = 2'b11;
			14'b00001000110011: M1r = 2'b11;
			14'b01001000110011: M1r = 2'b11;
			14'b10001000110011: M1r = 2'b11;
			14'b11001000110011: M1r = 2'b11;
			14'b00011000110011: M1r = 2'b11;
			14'b01011000110011: M1r = 2'b11;
			14'b10011000110011: M1r = 2'b11;
			14'b11011000110011: M1r = 2'b11;
			14'b00101000110011: M1r = 2'b11;
			14'b01101000110011: M1r = 2'b11;
			14'b10101000110011: M1r = 2'b11;
			14'b11101000110011: M1r = 2'b11;
			14'b00111000110011: M1r = 2'b11;
			14'b01111000110011: M1r = 2'b11;
			14'b10111000110011: M1r = 2'b11;
			14'b11111000110011: M1r = 2'b11;
			14'b00001100110011: M1r = 2'b11;
			14'b01001100110011: M1r = 2'b11;
			14'b10001100110011: M1r = 2'b11;
			14'b11001100110011: M1r = 2'b11;
			14'b00011100110011: M1r = 2'b11;
			14'b01011100110011: M1r = 2'b11;
			14'b10011100110011: M1r = 2'b11;
			14'b11011100110011: M1r = 2'b11;
			14'b00101100110011: M1r = 2'b11;
			14'b01101100110011: M1r = 2'b11;
			14'b10101100110011: M1r = 2'b11;
			14'b11101100110011: M1r = 2'b11;
			14'b00111100110011: M1r = 2'b11;
			14'b01111100110011: M1r = 2'b11;
			14'b10111100110011: M1r = 2'b11;
			14'b11111100110011: M1r = 2'b11;
			14'b00000001110011: M1r = 2'b11;
			14'b01000001110011: M1r = 2'b11;
			14'b10000001110011: M1r = 2'b11;
			14'b11000001110011: M1r = 2'b11;
			14'b00010001110011: M1r = 2'b11;
			14'b01010001110011: M1r = 2'b11;
			14'b10010001110011: M1r = 2'b11;
			14'b11010001110011: M1r = 2'b11;
			14'b00100001110011: M1r = 2'b10;
			14'b01100001110011: M1r = 2'b10;
			14'b10100001110011: M1r = 2'b10;
			14'b11100001110011: M1r = 2'b11;
			14'b00110001110011: M1r = 2'b10;
			14'b01110001110011: M1r = 2'b10;
			14'b10110001110011: M1r = 2'b10;
			14'b11110001110011: M1r = 2'b10;
			14'b00000101110011: M1r = 2'b11;
			14'b01000101110011: M1r = 2'b11;
			14'b10000101110011: M1r = 2'b11;
			14'b11000101110011: M1r = 2'b11;
			14'b00010101110011: M1r = 2'b11;
			14'b01010101110011: M1r = 2'b11;
			14'b10010101110011: M1r = 2'b11;
			14'b11010101110011: M1r = 2'b11;
			14'b00100101110011: M1r = 2'b11;
			14'b01100101110011: M1r = 2'b11;
			14'b10100101110011: M1r = 2'b11;
			14'b11100101110011: M1r = 2'b11;
			14'b00110101110011: M1r = 2'b10;
			14'b01110101110011: M1r = 2'b11;
			14'b10110101110011: M1r = 2'b11;
			14'b11110101110011: M1r = 2'b11;
			14'b00001001110011: M1r = 2'b11;
			14'b01001001110011: M1r = 2'b11;
			14'b10001001110011: M1r = 2'b11;
			14'b11001001110011: M1r = 2'b11;
			14'b00011001110011: M1r = 2'b11;
			14'b01011001110011: M1r = 2'b11;
			14'b10011001110011: M1r = 2'b11;
			14'b11011001110011: M1r = 2'b11;
			14'b00101001110011: M1r = 2'b11;
			14'b01101001110011: M1r = 2'b11;
			14'b10101001110011: M1r = 2'b11;
			14'b11101001110011: M1r = 2'b11;
			14'b00111001110011: M1r = 2'b11;
			14'b01111001110011: M1r = 2'b11;
			14'b10111001110011: M1r = 2'b11;
			14'b11111001110011: M1r = 2'b11;
			14'b00001101110011: M1r = 2'b11;
			14'b01001101110011: M1r = 2'b11;
			14'b10001101110011: M1r = 2'b11;
			14'b11001101110011: M1r = 2'b11;
			14'b00011101110011: M1r = 2'b11;
			14'b01011101110011: M1r = 2'b11;
			14'b10011101110011: M1r = 2'b11;
			14'b11011101110011: M1r = 2'b11;
			14'b00101101110011: M1r = 2'b11;
			14'b01101101110011: M1r = 2'b11;
			14'b10101101110011: M1r = 2'b11;
			14'b11101101110011: M1r = 2'b11;
			14'b00111101110011: M1r = 2'b11;
			14'b01111101110011: M1r = 2'b11;
			14'b10111101110011: M1r = 2'b11;
			14'b11111101110011: M1r = 2'b11;
			14'b00000010110011: M1r = 2'b11;
			14'b01000010110011: M1r = 2'b11;
			14'b10000010110011: M1r = 2'b11;
			14'b11000010110011: M1r = 2'b11;
			14'b00010010110011: M1r = 2'b10;
			14'b01010010110011: M1r = 2'b10;
			14'b10010010110011: M1r = 2'b11;
			14'b11010010110011: M1r = 2'b11;
			14'b00100010110011: M1r = 2'b10;
			14'b01100010110011: M1r = 2'b10;
			14'b10100010110011: M1r = 2'b10;
			14'b11100010110011: M1r = 2'b10;
			14'b00110010110011: M1r = 2'b01;
			14'b01110010110011: M1r = 2'b10;
			14'b10110010110011: M1r = 2'b10;
			14'b11110010110011: M1r = 2'b10;
			14'b00000110110011: M1r = 2'b11;
			14'b01000110110011: M1r = 2'b11;
			14'b10000110110011: M1r = 2'b11;
			14'b11000110110011: M1r = 2'b11;
			14'b00010110110011: M1r = 2'b11;
			14'b01010110110011: M1r = 2'b11;
			14'b10010110110011: M1r = 2'b11;
			14'b11010110110011: M1r = 2'b11;
			14'b00100110110011: M1r = 2'b11;
			14'b01100110110011: M1r = 2'b11;
			14'b10100110110011: M1r = 2'b11;
			14'b11100110110011: M1r = 2'b11;
			14'b00110110110011: M1r = 2'b10;
			14'b01110110110011: M1r = 2'b10;
			14'b10110110110011: M1r = 2'b10;
			14'b11110110110011: M1r = 2'b11;
			14'b00001010110011: M1r = 2'b11;
			14'b01001010110011: M1r = 2'b11;
			14'b10001010110011: M1r = 2'b11;
			14'b11001010110011: M1r = 2'b11;
			14'b00011010110011: M1r = 2'b11;
			14'b01011010110011: M1r = 2'b11;
			14'b10011010110011: M1r = 2'b11;
			14'b11011010110011: M1r = 2'b11;
			14'b00101010110011: M1r = 2'b11;
			14'b01101010110011: M1r = 2'b11;
			14'b10101010110011: M1r = 2'b11;
			14'b11101010110011: M1r = 2'b11;
			14'b00111010110011: M1r = 2'b11;
			14'b01111010110011: M1r = 2'b11;
			14'b10111010110011: M1r = 2'b11;
			14'b11111010110011: M1r = 2'b11;
			14'b00001110110011: M1r = 2'b11;
			14'b01001110110011: M1r = 2'b11;
			14'b10001110110011: M1r = 2'b11;
			14'b11001110110011: M1r = 2'b11;
			14'b00011110110011: M1r = 2'b11;
			14'b01011110110011: M1r = 2'b11;
			14'b10011110110011: M1r = 2'b11;
			14'b11011110110011: M1r = 2'b11;
			14'b00101110110011: M1r = 2'b11;
			14'b01101110110011: M1r = 2'b11;
			14'b10101110110011: M1r = 2'b11;
			14'b11101110110011: M1r = 2'b11;
			14'b00111110110011: M1r = 2'b11;
			14'b01111110110011: M1r = 2'b11;
			14'b10111110110011: M1r = 2'b11;
			14'b11111110110011: M1r = 2'b11;
			14'b00000011110011: M1r = 2'b11;
			14'b01000011110011: M1r = 2'b11;
			14'b10000011110011: M1r = 2'b11;
			14'b11000011110011: M1r = 2'b11;
			14'b00010011110011: M1r = 2'b10;
			14'b01010011110011: M1r = 2'b10;
			14'b10010011110011: M1r = 2'b10;
			14'b11010011110011: M1r = 2'b11;
			14'b00100011110011: M1r = 2'b10;
			14'b01100011110011: M1r = 2'b10;
			14'b10100011110011: M1r = 2'b10;
			14'b11100011110011: M1r = 2'b10;
			14'b00110011110011: M1r = 2'b01;
			14'b01110011110011: M1r = 2'b01;
			14'b10110011110011: M1r = 2'b01;
			14'b11110011110011: M1r = 2'b10;
			14'b00000111110011: M1r = 2'b11;
			14'b01000111110011: M1r = 2'b11;
			14'b10000111110011: M1r = 2'b11;
			14'b11000111110011: M1r = 2'b11;
			14'b00010111110011: M1r = 2'b11;
			14'b01010111110011: M1r = 2'b11;
			14'b10010111110011: M1r = 2'b11;
			14'b11010111110011: M1r = 2'b11;
			14'b00100111110011: M1r = 2'b10;
			14'b01100111110011: M1r = 2'b10;
			14'b10100111110011: M1r = 2'b11;
			14'b11100111110011: M1r = 2'b11;
			14'b00110111110011: M1r = 2'b10;
			14'b01110111110011: M1r = 2'b10;
			14'b10110111110011: M1r = 2'b10;
			14'b11110111110011: M1r = 2'b10;
			14'b00001011110011: M1r = 2'b11;
			14'b01001011110011: M1r = 2'b11;
			14'b10001011110011: M1r = 2'b11;
			14'b11001011110011: M1r = 2'b11;
			14'b00011011110011: M1r = 2'b11;
			14'b01011011110011: M1r = 2'b11;
			14'b10011011110011: M1r = 2'b11;
			14'b11011011110011: M1r = 2'b11;
			14'b00101011110011: M1r = 2'b11;
			14'b01101011110011: M1r = 2'b11;
			14'b10101011110011: M1r = 2'b11;
			14'b11101011110011: M1r = 2'b11;
			14'b00111011110011: M1r = 2'b11;
			14'b01111011110011: M1r = 2'b11;
			14'b10111011110011: M1r = 2'b11;
			14'b11111011110011: M1r = 2'b11;
			14'b00001111110011: M1r = 2'b11;
			14'b01001111110011: M1r = 2'b11;
			14'b10001111110011: M1r = 2'b11;
			14'b11001111110011: M1r = 2'b11;
			14'b00011111110011: M1r = 2'b11;
			14'b01011111110011: M1r = 2'b11;
			14'b10011111110011: M1r = 2'b11;
			14'b11011111110011: M1r = 2'b11;
			14'b00101111110011: M1r = 2'b11;
			14'b01101111110011: M1r = 2'b11;
			14'b10101111110011: M1r = 2'b11;
			14'b11101111110011: M1r = 2'b11;
			14'b00111111110011: M1r = 2'b11;
			14'b01111111110011: M1r = 2'b11;
			14'b10111111110011: M1r = 2'b11;
			14'b11111111110011: M1r = 2'b11;
			14'b00000000000111: M1r = 2'b01;
			14'b01000000000111: M1r = 2'b01;
			14'b10000000000111: M1r = 2'b10;
			14'b11000000000111: M1r = 2'b10;
			14'b00010000000111: M1r = 2'b01;
			14'b01010000000111: M1r = 2'b01;
			14'b10010000000111: M1r = 2'b01;
			14'b11010000000111: M1r = 2'b01;
			14'b00100000000111: M1r = 2'b00;
			14'b01100000000111: M1r = 2'b00;
			14'b10100000000111: M1r = 2'b01;
			14'b11100000000111: M1r = 2'b01;
			14'b00110000000111: M1r = 2'b00;
			14'b01110000000111: M1r = 2'b00;
			14'b10110000000111: M1r = 2'b00;
			14'b11110000000111: M1r = 2'b00;
			14'b00000100000111: M1r = 2'b10;
			14'b01000100000111: M1r = 2'b10;
			14'b10000100000111: M1r = 2'b10;
			14'b11000100000111: M1r = 2'b10;
			14'b00010100000111: M1r = 2'b10;
			14'b01010100000111: M1r = 2'b10;
			14'b10010100000111: M1r = 2'b10;
			14'b11010100000111: M1r = 2'b10;
			14'b00100100000111: M1r = 2'b01;
			14'b01100100000111: M1r = 2'b01;
			14'b10100100000111: M1r = 2'b01;
			14'b11100100000111: M1r = 2'b10;
			14'b00110100000111: M1r = 2'b01;
			14'b01110100000111: M1r = 2'b01;
			14'b10110100000111: M1r = 2'b01;
			14'b11110100000111: M1r = 2'b01;
			14'b00001000000111: M1r = 2'b11;
			14'b01001000000111: M1r = 2'b11;
			14'b10001000000111: M1r = 2'b11;
			14'b11001000000111: M1r = 2'b11;
			14'b00011000000111: M1r = 2'b10;
			14'b01011000000111: M1r = 2'b10;
			14'b10011000000111: M1r = 2'b11;
			14'b11011000000111: M1r = 2'b11;
			14'b00101000000111: M1r = 2'b10;
			14'b01101000000111: M1r = 2'b10;
			14'b10101000000111: M1r = 2'b10;
			14'b11101000000111: M1r = 2'b10;
			14'b00111000000111: M1r = 2'b01;
			14'b01111000000111: M1r = 2'b01;
			14'b10111000000111: M1r = 2'b10;
			14'b11111000000111: M1r = 2'b10;
			14'b00001100000111: M1r = 2'b11;
			14'b01001100000111: M1r = 2'b11;
			14'b10001100000111: M1r = 2'b11;
			14'b11001100000111: M1r = 2'b11;
			14'b00011100000111: M1r = 2'b11;
			14'b01011100000111: M1r = 2'b11;
			14'b10011100000111: M1r = 2'b11;
			14'b11011100000111: M1r = 2'b11;
			14'b00101100000111: M1r = 2'b11;
			14'b01101100000111: M1r = 2'b11;
			14'b10101100000111: M1r = 2'b11;
			14'b11101100000111: M1r = 2'b11;
			14'b00111100000111: M1r = 2'b10;
			14'b01111100000111: M1r = 2'b10;
			14'b10111100000111: M1r = 2'b10;
			14'b11111100000111: M1r = 2'b11;
			14'b00000001000111: M1r = 2'b01;
			14'b01000001000111: M1r = 2'b01;
			14'b10000001000111: M1r = 2'b01;
			14'b11000001000111: M1r = 2'b01;
			14'b00010001000111: M1r = 2'b01;
			14'b01010001000111: M1r = 2'b01;
			14'b10010001000111: M1r = 2'b01;
			14'b11010001000111: M1r = 2'b01;
			14'b00100001000111: M1r = 2'b00;
			14'b01100001000111: M1r = 2'b00;
			14'b10100001000111: M1r = 2'b00;
			14'b11100001000111: M1r = 2'b01;
			14'b00110001000111: M1r = 2'b00;
			14'b01110001000111: M1r = 2'b00;
			14'b10110001000111: M1r = 2'b00;
			14'b11110001000111: M1r = 2'b00;
			14'b00000101000111: M1r = 2'b10;
			14'b01000101000111: M1r = 2'b10;
			14'b10000101000111: M1r = 2'b10;
			14'b11000101000111: M1r = 2'b10;
			14'b00010101000111: M1r = 2'b01;
			14'b01010101000111: M1r = 2'b01;
			14'b10010101000111: M1r = 2'b10;
			14'b11010101000111: M1r = 2'b10;
			14'b00100101000111: M1r = 2'b01;
			14'b01100101000111: M1r = 2'b01;
			14'b10100101000111: M1r = 2'b01;
			14'b11100101000111: M1r = 2'b01;
			14'b00110101000111: M1r = 2'b00;
			14'b01110101000111: M1r = 2'b00;
			14'b10110101000111: M1r = 2'b01;
			14'b11110101000111: M1r = 2'b01;
			14'b00001001000111: M1r = 2'b10;
			14'b01001001000111: M1r = 2'b11;
			14'b10001001000111: M1r = 2'b11;
			14'b11001001000111: M1r = 2'b11;
			14'b00011001000111: M1r = 2'b10;
			14'b01011001000111: M1r = 2'b10;
			14'b10011001000111: M1r = 2'b10;
			14'b11011001000111: M1r = 2'b10;
			14'b00101001000111: M1r = 2'b10;
			14'b01101001000111: M1r = 2'b10;
			14'b10101001000111: M1r = 2'b10;
			14'b11101001000111: M1r = 2'b10;
			14'b00111001000111: M1r = 2'b01;
			14'b01111001000111: M1r = 2'b01;
			14'b10111001000111: M1r = 2'b01;
			14'b11111001000111: M1r = 2'b10;
			14'b00001101000111: M1r = 2'b11;
			14'b01001101000111: M1r = 2'b11;
			14'b10001101000111: M1r = 2'b11;
			14'b11001101000111: M1r = 2'b11;
			14'b00011101000111: M1r = 2'b11;
			14'b01011101000111: M1r = 2'b11;
			14'b10011101000111: M1r = 2'b11;
			14'b11011101000111: M1r = 2'b11;
			14'b00101101000111: M1r = 2'b10;
			14'b01101101000111: M1r = 2'b10;
			14'b10101101000111: M1r = 2'b11;
			14'b11101101000111: M1r = 2'b11;
			14'b00111101000111: M1r = 2'b10;
			14'b01111101000111: M1r = 2'b10;
			14'b10111101000111: M1r = 2'b10;
			14'b11111101000111: M1r = 2'b10;
			14'b00000010000111: M1r = 2'b01;
			14'b01000010000111: M1r = 2'b01;
			14'b10000010000111: M1r = 2'b01;
			14'b11000010000111: M1r = 2'b01;
			14'b00010010000111: M1r = 2'b00;
			14'b01010010000111: M1r = 2'b00;
			14'b10010010000111: M1r = 2'b01;
			14'b11010010000111: M1r = 2'b01;
			14'b00100010000111: M1r = 2'b00;
			14'b01100010000111: M1r = 2'b00;
			14'b10100010000111: M1r = 2'b00;
			14'b11100010000111: M1r = 2'b00;
			14'b00110010000111: M1r = 2'b00;
			14'b01110010000111: M1r = 2'b00;
			14'b10110010000111: M1r = 2'b00;
			14'b11110010000111: M1r = 2'b00;
			14'b00000110000111: M1r = 2'b01;
			14'b01000110000111: M1r = 2'b10;
			14'b10000110000111: M1r = 2'b10;
			14'b11000110000111: M1r = 2'b10;
			14'b00010110000111: M1r = 2'b01;
			14'b01010110000111: M1r = 2'b01;
			14'b10010110000111: M1r = 2'b01;
			14'b11010110000111: M1r = 2'b01;
			14'b00100110000111: M1r = 2'b01;
			14'b01100110000111: M1r = 2'b01;
			14'b10100110000111: M1r = 2'b01;
			14'b11100110000111: M1r = 2'b01;
			14'b00110110000111: M1r = 2'b00;
			14'b01110110000111: M1r = 2'b00;
			14'b10110110000111: M1r = 2'b00;
			14'b11110110000111: M1r = 2'b01;
			14'b00001010000111: M1r = 2'b10;
			14'b01001010000111: M1r = 2'b10;
			14'b10001010000111: M1r = 2'b11;
			14'b11001010000111: M1r = 2'b11;
			14'b00011010000111: M1r = 2'b10;
			14'b01011010000111: M1r = 2'b10;
			14'b10011010000111: M1r = 2'b10;
			14'b11011010000111: M1r = 2'b10;
			14'b00101010000111: M1r = 2'b01;
			14'b01101010000111: M1r = 2'b01;
			14'b10101010000111: M1r = 2'b10;
			14'b11101010000111: M1r = 2'b10;
			14'b00111010000111: M1r = 2'b01;
			14'b01111010000111: M1r = 2'b01;
			14'b10111010000111: M1r = 2'b01;
			14'b11111010000111: M1r = 2'b01;
			14'b00001110000111: M1r = 2'b11;
			14'b01001110000111: M1r = 2'b11;
			14'b10001110000111: M1r = 2'b11;
			14'b11001110000111: M1r = 2'b11;
			14'b00011110000111: M1r = 2'b10;
			14'b01011110000111: M1r = 2'b11;
			14'b10011110000111: M1r = 2'b11;
			14'b11011110000111: M1r = 2'b11;
			14'b00101110000111: M1r = 2'b10;
			14'b01101110000111: M1r = 2'b10;
			14'b10101110000111: M1r = 2'b10;
			14'b11101110000111: M1r = 2'b10;
			14'b00111110000111: M1r = 2'b10;
			14'b01111110000111: M1r = 2'b10;
			14'b10111110000111: M1r = 2'b10;
			14'b11111110000111: M1r = 2'b10;
			14'b00000011000111: M1r = 2'b00;
			14'b01000011000111: M1r = 2'b01;
			14'b10000011000111: M1r = 2'b01;
			14'b11000011000111: M1r = 2'b01;
			14'b00010011000111: M1r = 2'b00;
			14'b01010011000111: M1r = 2'b00;
			14'b10010011000111: M1r = 2'b00;
			14'b11010011000111: M1r = 2'b00;
			14'b00100011000111: M1r = 2'b00;
			14'b01100011000111: M1r = 2'b00;
			14'b10100011000111: M1r = 2'b00;
			14'b11100011000111: M1r = 2'b00;
			14'b00110011000111: M1r = 2'b00;
			14'b01110011000111: M1r = 2'b00;
			14'b10110011000111: M1r = 2'b00;
			14'b11110011000111: M1r = 2'b00;
			14'b00000111000111: M1r = 2'b01;
			14'b01000111000111: M1r = 2'b01;
			14'b10000111000111: M1r = 2'b01;
			14'b11000111000111: M1r = 2'b10;
			14'b00010111000111: M1r = 2'b01;
			14'b01010111000111: M1r = 2'b01;
			14'b10010111000111: M1r = 2'b01;
			14'b11010111000111: M1r = 2'b01;
			14'b00100111000111: M1r = 2'b00;
			14'b01100111000111: M1r = 2'b00;
			14'b10100111000111: M1r = 2'b01;
			14'b11100111000111: M1r = 2'b01;
			14'b00110111000111: M1r = 2'b00;
			14'b01110111000111: M1r = 2'b00;
			14'b10110111000111: M1r = 2'b00;
			14'b11110111000111: M1r = 2'b00;
			14'b00001011000111: M1r = 2'b10;
			14'b01001011000111: M1r = 2'b10;
			14'b10001011000111: M1r = 2'b10;
			14'b11001011000111: M1r = 2'b10;
			14'b00011011000111: M1r = 2'b01;
			14'b01011011000111: M1r = 2'b10;
			14'b10011011000111: M1r = 2'b10;
			14'b11011011000111: M1r = 2'b10;
			14'b00101011000111: M1r = 2'b01;
			14'b01101011000111: M1r = 2'b01;
			14'b10101011000111: M1r = 2'b01;
			14'b11101011000111: M1r = 2'b01;
			14'b00111011000111: M1r = 2'b01;
			14'b01111011000111: M1r = 2'b01;
			14'b10111011000111: M1r = 2'b01;
			14'b11111011000111: M1r = 2'b01;
			14'b00001111000111: M1r = 2'b11;
			14'b01001111000111: M1r = 2'b11;
			14'b10001111000111: M1r = 2'b11;
			14'b11001111000111: M1r = 2'b11;
			14'b00011111000111: M1r = 2'b10;
			14'b01011111000111: M1r = 2'b10;
			14'b10011111000111: M1r = 2'b11;
			14'b11011111000111: M1r = 2'b11;
			14'b00101111000111: M1r = 2'b10;
			14'b01101111000111: M1r = 2'b10;
			14'b10101111000111: M1r = 2'b10;
			14'b11101111000111: M1r = 2'b10;
			14'b00111111000111: M1r = 2'b01;
			14'b01111111000111: M1r = 2'b01;
			14'b10111111000111: M1r = 2'b10;
			14'b11111111000111: M1r = 2'b10;
			14'b00000000010111: M1r = 2'b10;
			14'b01000000010111: M1r = 2'b10;
			14'b10000000010111: M1r = 2'b10;
			14'b11000000010111: M1r = 2'b10;
			14'b00010000010111: M1r = 2'b01;
			14'b01010000010111: M1r = 2'b01;
			14'b10010000010111: M1r = 2'b10;
			14'b11010000010111: M1r = 2'b10;
			14'b00100000010111: M1r = 2'b01;
			14'b01100000010111: M1r = 2'b01;
			14'b10100000010111: M1r = 2'b01;
			14'b11100000010111: M1r = 2'b01;
			14'b00110000010111: M1r = 2'b00;
			14'b01110000010111: M1r = 2'b00;
			14'b10110000010111: M1r = 2'b01;
			14'b11110000010111: M1r = 2'b01;
			14'b00000100010111: M1r = 2'b10;
			14'b01000100010111: M1r = 2'b11;
			14'b10000100010111: M1r = 2'b11;
			14'b11000100010111: M1r = 2'b11;
			14'b00010100010111: M1r = 2'b10;
			14'b01010100010111: M1r = 2'b10;
			14'b10010100010111: M1r = 2'b10;
			14'b11010100010111: M1r = 2'b10;
			14'b00100100010111: M1r = 2'b10;
			14'b01100100010111: M1r = 2'b10;
			14'b10100100010111: M1r = 2'b10;
			14'b11100100010111: M1r = 2'b10;
			14'b00110100010111: M1r = 2'b01;
			14'b01110100010111: M1r = 2'b01;
			14'b10110100010111: M1r = 2'b01;
			14'b11110100010111: M1r = 2'b01;
			14'b00001000010111: M1r = 2'b11;
			14'b01001000010111: M1r = 2'b11;
			14'b10001000010111: M1r = 2'b11;
			14'b11001000010111: M1r = 2'b11;
			14'b00011000010111: M1r = 2'b11;
			14'b01011000010111: M1r = 2'b11;
			14'b10011000010111: M1r = 2'b11;
			14'b11011000010111: M1r = 2'b11;
			14'b00101000010111: M1r = 2'b10;
			14'b01101000010111: M1r = 2'b10;
			14'b10101000010111: M1r = 2'b11;
			14'b11101000010111: M1r = 2'b11;
			14'b00111000010111: M1r = 2'b10;
			14'b01111000010111: M1r = 2'b10;
			14'b10111000010111: M1r = 2'b10;
			14'b11111000010111: M1r = 2'b10;
			14'b00001100010111: M1r = 2'b11;
			14'b01001100010111: M1r = 2'b11;
			14'b10001100010111: M1r = 2'b11;
			14'b11001100010111: M1r = 2'b11;
			14'b00011100010111: M1r = 2'b11;
			14'b01011100010111: M1r = 2'b11;
			14'b10011100010111: M1r = 2'b11;
			14'b11011100010111: M1r = 2'b11;
			14'b00101100010111: M1r = 2'b11;
			14'b01101100010111: M1r = 2'b11;
			14'b10101100010111: M1r = 2'b11;
			14'b11101100010111: M1r = 2'b11;
			14'b00111100010111: M1r = 2'b11;
			14'b01111100010111: M1r = 2'b11;
			14'b10111100010111: M1r = 2'b11;
			14'b11111100010111: M1r = 2'b11;
			14'b00000001010111: M1r = 2'b01;
			14'b01000001010111: M1r = 2'b10;
			14'b10000001010111: M1r = 2'b10;
			14'b11000001010111: M1r = 2'b10;
			14'b00010001010111: M1r = 2'b01;
			14'b01010001010111: M1r = 2'b01;
			14'b10010001010111: M1r = 2'b01;
			14'b11010001010111: M1r = 2'b01;
			14'b00100001010111: M1r = 2'b00;
			14'b01100001010111: M1r = 2'b01;
			14'b10100001010111: M1r = 2'b01;
			14'b11100001010111: M1r = 2'b01;
			14'b00110001010111: M1r = 2'b00;
			14'b01110001010111: M1r = 2'b00;
			14'b10110001010111: M1r = 2'b00;
			14'b11110001010111: M1r = 2'b00;
			14'b00000101010111: M1r = 2'b10;
			14'b01000101010111: M1r = 2'b10;
			14'b10000101010111: M1r = 2'b10;
			14'b11000101010111: M1r = 2'b11;
			14'b00010101010111: M1r = 2'b10;
			14'b01010101010111: M1r = 2'b10;
			14'b10010101010111: M1r = 2'b10;
			14'b11010101010111: M1r = 2'b10;
			14'b00100101010111: M1r = 2'b01;
			14'b01100101010111: M1r = 2'b01;
			14'b10100101010111: M1r = 2'b10;
			14'b11100101010111: M1r = 2'b10;
			14'b00110101010111: M1r = 2'b01;
			14'b01110101010111: M1r = 2'b01;
			14'b10110101010111: M1r = 2'b01;
			14'b11110101010111: M1r = 2'b01;
			14'b00001001010111: M1r = 2'b11;
			14'b01001001010111: M1r = 2'b11;
			14'b10001001010111: M1r = 2'b11;
			14'b11001001010111: M1r = 2'b11;
			14'b00011001010111: M1r = 2'b10;
			14'b01011001010111: M1r = 2'b11;
			14'b10011001010111: M1r = 2'b11;
			14'b11011001010111: M1r = 2'b11;
			14'b00101001010111: M1r = 2'b10;
			14'b01101001010111: M1r = 2'b10;
			14'b10101001010111: M1r = 2'b10;
			14'b11101001010111: M1r = 2'b10;
			14'b00111001010111: M1r = 2'b10;
			14'b01111001010111: M1r = 2'b10;
			14'b10111001010111: M1r = 2'b10;
			14'b11111001010111: M1r = 2'b10;
			14'b00001101010111: M1r = 2'b11;
			14'b01001101010111: M1r = 2'b11;
			14'b10001101010111: M1r = 2'b11;
			14'b11001101010111: M1r = 2'b11;
			14'b00011101010111: M1r = 2'b11;
			14'b01011101010111: M1r = 2'b11;
			14'b10011101010111: M1r = 2'b11;
			14'b11011101010111: M1r = 2'b11;
			14'b00101101010111: M1r = 2'b11;
			14'b01101101010111: M1r = 2'b11;
			14'b10101101010111: M1r = 2'b11;
			14'b11101101010111: M1r = 2'b11;
			14'b00111101010111: M1r = 2'b10;
			14'b01111101010111: M1r = 2'b10;
			14'b10111101010111: M1r = 2'b11;
			14'b11111101010111: M1r = 2'b11;
			14'b00000010010111: M1r = 2'b01;
			14'b01000010010111: M1r = 2'b01;
			14'b10000010010111: M1r = 2'b01;
			14'b11000010010111: M1r = 2'b10;
			14'b00010010010111: M1r = 2'b01;
			14'b01010010010111: M1r = 2'b01;
			14'b10010010010111: M1r = 2'b01;
			14'b11010010010111: M1r = 2'b01;
			14'b00100010010111: M1r = 2'b00;
			14'b01100010010111: M1r = 2'b00;
			14'b10100010010111: M1r = 2'b01;
			14'b11100010010111: M1r = 2'b01;
			14'b00110010010111: M1r = 2'b00;
			14'b01110010010111: M1r = 2'b00;
			14'b10110010010111: M1r = 2'b00;
			14'b11110010010111: M1r = 2'b00;
			14'b00000110010111: M1r = 2'b10;
			14'b01000110010111: M1r = 2'b10;
			14'b10000110010111: M1r = 2'b10;
			14'b11000110010111: M1r = 2'b10;
			14'b00010110010111: M1r = 2'b01;
			14'b01010110010111: M1r = 2'b10;
			14'b10010110010111: M1r = 2'b10;
			14'b11010110010111: M1r = 2'b10;
			14'b00100110010111: M1r = 2'b01;
			14'b01100110010111: M1r = 2'b01;
			14'b10100110010111: M1r = 2'b01;
			14'b11100110010111: M1r = 2'b01;
			14'b00110110010111: M1r = 2'b00;
			14'b01110110010111: M1r = 2'b01;
			14'b10110110010111: M1r = 2'b01;
			14'b11110110010111: M1r = 2'b01;
			14'b00001010010111: M1r = 2'b11;
			14'b01001010010111: M1r = 2'b11;
			14'b10001010010111: M1r = 2'b11;
			14'b11001010010111: M1r = 2'b11;
			14'b00011010010111: M1r = 2'b10;
			14'b01011010010111: M1r = 2'b10;
			14'b10011010010111: M1r = 2'b10;
			14'b11011010010111: M1r = 2'b11;
			14'b00101010010111: M1r = 2'b10;
			14'b01101010010111: M1r = 2'b10;
			14'b10101010010111: M1r = 2'b10;
			14'b11101010010111: M1r = 2'b10;
			14'b00111010010111: M1r = 2'b01;
			14'b01111010010111: M1r = 2'b01;
			14'b10111010010111: M1r = 2'b10;
			14'b11111010010111: M1r = 2'b10;
			14'b00001110010111: M1r = 2'b11;
			14'b01001110010111: M1r = 2'b11;
			14'b10001110010111: M1r = 2'b11;
			14'b11001110010111: M1r = 2'b11;
			14'b00011110010111: M1r = 2'b11;
			14'b01011110010111: M1r = 2'b11;
			14'b10011110010111: M1r = 2'b11;
			14'b11011110010111: M1r = 2'b11;
			14'b00101110010111: M1r = 2'b10;
			14'b01101110010111: M1r = 2'b11;
			14'b10101110010111: M1r = 2'b11;
			14'b11101110010111: M1r = 2'b11;
			14'b00111110010111: M1r = 2'b10;
			14'b01111110010111: M1r = 2'b10;
			14'b10111110010111: M1r = 2'b10;
			14'b11111110010111: M1r = 2'b10;
			14'b00000011010111: M1r = 2'b01;
			14'b01000011010111: M1r = 2'b01;
			14'b10000011010111: M1r = 2'b01;
			14'b11000011010111: M1r = 2'b01;
			14'b00010011010111: M1r = 2'b00;
			14'b01010011010111: M1r = 2'b01;
			14'b10010011010111: M1r = 2'b01;
			14'b11010011010111: M1r = 2'b01;
			14'b00100011010111: M1r = 2'b00;
			14'b01100011010111: M1r = 2'b00;
			14'b10100011010111: M1r = 2'b00;
			14'b11100011010111: M1r = 2'b00;
			14'b00110011010111: M1r = 2'b00;
			14'b01110011010111: M1r = 2'b00;
			14'b10110011010111: M1r = 2'b00;
			14'b11110011010111: M1r = 2'b00;
			14'b00000111010111: M1r = 2'b10;
			14'b01000111010111: M1r = 2'b10;
			14'b10000111010111: M1r = 2'b10;
			14'b11000111010111: M1r = 2'b10;
			14'b00010111010111: M1r = 2'b01;
			14'b01010111010111: M1r = 2'b01;
			14'b10010111010111: M1r = 2'b01;
			14'b11010111010111: M1r = 2'b10;
			14'b00100111010111: M1r = 2'b01;
			14'b01100111010111: M1r = 2'b01;
			14'b10100111010111: M1r = 2'b01;
			14'b11100111010111: M1r = 2'b01;
			14'b00110111010111: M1r = 2'b00;
			14'b01110111010111: M1r = 2'b00;
			14'b10110111010111: M1r = 2'b01;
			14'b11110111010111: M1r = 2'b01;
			14'b00001011010111: M1r = 2'b10;
			14'b01001011010111: M1r = 2'b11;
			14'b10001011010111: M1r = 2'b11;
			14'b11001011010111: M1r = 2'b11;
			14'b00011011010111: M1r = 2'b10;
			14'b01011011010111: M1r = 2'b10;
			14'b10011011010111: M1r = 2'b10;
			14'b11011011010111: M1r = 2'b10;
			14'b00101011010111: M1r = 2'b01;
			14'b01101011010111: M1r = 2'b10;
			14'b10101011010111: M1r = 2'b10;
			14'b11101011010111: M1r = 2'b10;
			14'b00111011010111: M1r = 2'b01;
			14'b01111011010111: M1r = 2'b01;
			14'b10111011010111: M1r = 2'b01;
			14'b11111011010111: M1r = 2'b01;
			14'b00001111010111: M1r = 2'b11;
			14'b01001111010111: M1r = 2'b11;
			14'b10001111010111: M1r = 2'b11;
			14'b11001111010111: M1r = 2'b11;
			14'b00011111010111: M1r = 2'b11;
			14'b01011111010111: M1r = 2'b11;
			14'b10011111010111: M1r = 2'b11;
			14'b11011111010111: M1r = 2'b11;
			14'b00101111010111: M1r = 2'b10;
			14'b01101111010111: M1r = 2'b10;
			14'b10101111010111: M1r = 2'b10;
			14'b11101111010111: M1r = 2'b11;
			14'b00111111010111: M1r = 2'b10;
			14'b01111111010111: M1r = 2'b10;
			14'b10111111010111: M1r = 2'b10;
			14'b11111111010111: M1r = 2'b10;
			14'b00000000100111: M1r = 2'b10;
			14'b01000000100111: M1r = 2'b10;
			14'b10000000100111: M1r = 2'b10;
			14'b11000000100111: M1r = 2'b11;
			14'b00010000100111: M1r = 2'b10;
			14'b01010000100111: M1r = 2'b10;
			14'b10010000100111: M1r = 2'b10;
			14'b11010000100111: M1r = 2'b10;
			14'b00100000100111: M1r = 2'b01;
			14'b01100000100111: M1r = 2'b01;
			14'b10100000100111: M1r = 2'b01;
			14'b11100000100111: M1r = 2'b10;
			14'b00110000100111: M1r = 2'b01;
			14'b01110000100111: M1r = 2'b01;
			14'b10110000100111: M1r = 2'b01;
			14'b11110000100111: M1r = 2'b01;
			14'b00000100100111: M1r = 2'b11;
			14'b01000100100111: M1r = 2'b11;
			14'b10000100100111: M1r = 2'b11;
			14'b11000100100111: M1r = 2'b11;
			14'b00010100100111: M1r = 2'b10;
			14'b01010100100111: M1r = 2'b11;
			14'b10010100100111: M1r = 2'b11;
			14'b11010100100111: M1r = 2'b11;
			14'b00100100100111: M1r = 2'b10;
			14'b01100100100111: M1r = 2'b10;
			14'b10100100100111: M1r = 2'b10;
			14'b11100100100111: M1r = 2'b10;
			14'b00110100100111: M1r = 2'b01;
			14'b01110100100111: M1r = 2'b10;
			14'b10110100100111: M1r = 2'b10;
			14'b11110100100111: M1r = 2'b10;
			14'b00001000100111: M1r = 2'b11;
			14'b01001000100111: M1r = 2'b11;
			14'b10001000100111: M1r = 2'b11;
			14'b11001000100111: M1r = 2'b11;
			14'b00011000100111: M1r = 2'b11;
			14'b01011000100111: M1r = 2'b11;
			14'b10011000100111: M1r = 2'b11;
			14'b11011000100111: M1r = 2'b11;
			14'b00101000100111: M1r = 2'b11;
			14'b01101000100111: M1r = 2'b11;
			14'b10101000100111: M1r = 2'b11;
			14'b11101000100111: M1r = 2'b11;
			14'b00111000100111: M1r = 2'b10;
			14'b01111000100111: M1r = 2'b10;
			14'b10111000100111: M1r = 2'b11;
			14'b11111000100111: M1r = 2'b11;
			14'b00001100100111: M1r = 2'b11;
			14'b01001100100111: M1r = 2'b11;
			14'b10001100100111: M1r = 2'b11;
			14'b11001100100111: M1r = 2'b11;
			14'b00011100100111: M1r = 2'b11;
			14'b01011100100111: M1r = 2'b11;
			14'b10011100100111: M1r = 2'b11;
			14'b11011100100111: M1r = 2'b11;
			14'b00101100100111: M1r = 2'b11;
			14'b01101100100111: M1r = 2'b11;
			14'b10101100100111: M1r = 2'b11;
			14'b11101100100111: M1r = 2'b11;
			14'b00111100100111: M1r = 2'b11;
			14'b01111100100111: M1r = 2'b11;
			14'b10111100100111: M1r = 2'b11;
			14'b11111100100111: M1r = 2'b11;
			14'b00000001100111: M1r = 2'b10;
			14'b01000001100111: M1r = 2'b10;
			14'b10000001100111: M1r = 2'b10;
			14'b11000001100111: M1r = 2'b10;
			14'b00010001100111: M1r = 2'b01;
			14'b01010001100111: M1r = 2'b10;
			14'b10010001100111: M1r = 2'b10;
			14'b11010001100111: M1r = 2'b10;
			14'b00100001100111: M1r = 2'b01;
			14'b01100001100111: M1r = 2'b01;
			14'b10100001100111: M1r = 2'b01;
			14'b11100001100111: M1r = 2'b01;
			14'b00110001100111: M1r = 2'b00;
			14'b01110001100111: M1r = 2'b01;
			14'b10110001100111: M1r = 2'b01;
			14'b11110001100111: M1r = 2'b01;
			14'b00000101100111: M1r = 2'b11;
			14'b01000101100111: M1r = 2'b11;
			14'b10000101100111: M1r = 2'b11;
			14'b11000101100111: M1r = 2'b11;
			14'b00010101100111: M1r = 2'b10;
			14'b01010101100111: M1r = 2'b10;
			14'b10010101100111: M1r = 2'b10;
			14'b11010101100111: M1r = 2'b11;
			14'b00100101100111: M1r = 2'b10;
			14'b01100101100111: M1r = 2'b10;
			14'b10100101100111: M1r = 2'b10;
			14'b11100101100111: M1r = 2'b10;
			14'b00110101100111: M1r = 2'b01;
			14'b01110101100111: M1r = 2'b01;
			14'b10110101100111: M1r = 2'b01;
			14'b11110101100111: M1r = 2'b10;
			14'b00001001100111: M1r = 2'b11;
			14'b01001001100111: M1r = 2'b11;
			14'b10001001100111: M1r = 2'b11;
			14'b11001001100111: M1r = 2'b11;
			14'b00011001100111: M1r = 2'b11;
			14'b01011001100111: M1r = 2'b11;
			14'b10011001100111: M1r = 2'b11;
			14'b11011001100111: M1r = 2'b11;
			14'b00101001100111: M1r = 2'b10;
			14'b01101001100111: M1r = 2'b11;
			14'b10101001100111: M1r = 2'b11;
			14'b11101001100111: M1r = 2'b11;
			14'b00111001100111: M1r = 2'b10;
			14'b01111001100111: M1r = 2'b10;
			14'b10111001100111: M1r = 2'b10;
			14'b11111001100111: M1r = 2'b10;
			14'b00001101100111: M1r = 2'b11;
			14'b01001101100111: M1r = 2'b11;
			14'b10001101100111: M1r = 2'b11;
			14'b11001101100111: M1r = 2'b11;
			14'b00011101100111: M1r = 2'b11;
			14'b01011101100111: M1r = 2'b11;
			14'b10011101100111: M1r = 2'b11;
			14'b11011101100111: M1r = 2'b11;
			14'b00101101100111: M1r = 2'b11;
			14'b01101101100111: M1r = 2'b11;
			14'b10101101100111: M1r = 2'b11;
			14'b11101101100111: M1r = 2'b11;
			14'b00111101100111: M1r = 2'b11;
			14'b01111101100111: M1r = 2'b11;
			14'b10111101100111: M1r = 2'b11;
			14'b11111101100111: M1r = 2'b11;
			14'b00000010100111: M1r = 2'b10;
			14'b01000010100111: M1r = 2'b10;
			14'b10000010100111: M1r = 2'b10;
			14'b11000010100111: M1r = 2'b10;
			14'b00010010100111: M1r = 2'b01;
			14'b01010010100111: M1r = 2'b01;
			14'b10010010100111: M1r = 2'b01;
			14'b11010010100111: M1r = 2'b10;
			14'b00100010100111: M1r = 2'b01;
			14'b01100010100111: M1r = 2'b01;
			14'b10100010100111: M1r = 2'b01;
			14'b11100010100111: M1r = 2'b01;
			14'b00110010100111: M1r = 2'b00;
			14'b01110010100111: M1r = 2'b00;
			14'b10110010100111: M1r = 2'b00;
			14'b11110010100111: M1r = 2'b01;
			14'b00000110100111: M1r = 2'b10;
			14'b01000110100111: M1r = 2'b10;
			14'b10000110100111: M1r = 2'b11;
			14'b11000110100111: M1r = 2'b11;
			14'b00010110100111: M1r = 2'b10;
			14'b01010110100111: M1r = 2'b10;
			14'b10010110100111: M1r = 2'b10;
			14'b11010110100111: M1r = 2'b10;
			14'b00100110100111: M1r = 2'b01;
			14'b01100110100111: M1r = 2'b10;
			14'b10100110100111: M1r = 2'b10;
			14'b11100110100111: M1r = 2'b10;
			14'b00110110100111: M1r = 2'b01;
			14'b01110110100111: M1r = 2'b01;
			14'b10110110100111: M1r = 2'b01;
			14'b11110110100111: M1r = 2'b01;
			14'b00001010100111: M1r = 2'b11;
			14'b01001010100111: M1r = 2'b11;
			14'b10001010100111: M1r = 2'b11;
			14'b11001010100111: M1r = 2'b11;
			14'b00011010100111: M1r = 2'b11;
			14'b01011010100111: M1r = 2'b11;
			14'b10011010100111: M1r = 2'b11;
			14'b11011010100111: M1r = 2'b11;
			14'b00101010100111: M1r = 2'b10;
			14'b01101010100111: M1r = 2'b10;
			14'b10101010100111: M1r = 2'b10;
			14'b11101010100111: M1r = 2'b11;
			14'b00111010100111: M1r = 2'b10;
			14'b01111010100111: M1r = 2'b10;
			14'b10111010100111: M1r = 2'b10;
			14'b11111010100111: M1r = 2'b10;
			14'b00001110100111: M1r = 2'b11;
			14'b01001110100111: M1r = 2'b11;
			14'b10001110100111: M1r = 2'b11;
			14'b11001110100111: M1r = 2'b11;
			14'b00011110100111: M1r = 2'b11;
			14'b01011110100111: M1r = 2'b11;
			14'b10011110100111: M1r = 2'b11;
			14'b11011110100111: M1r = 2'b11;
			14'b00101110100111: M1r = 2'b11;
			14'b01101110100111: M1r = 2'b11;
			14'b10101110100111: M1r = 2'b11;
			14'b11101110100111: M1r = 2'b11;
			14'b00111110100111: M1r = 2'b10;
			14'b01111110100111: M1r = 2'b11;
			14'b10111110100111: M1r = 2'b11;
			14'b11111110100111: M1r = 2'b11;
			14'b00000011100111: M1r = 2'b01;
			14'b01000011100111: M1r = 2'b01;
			14'b10000011100111: M1r = 2'b10;
			14'b11000011100111: M1r = 2'b10;
			14'b00010011100111: M1r = 2'b01;
			14'b01010011100111: M1r = 2'b01;
			14'b10010011100111: M1r = 2'b01;
			14'b11010011100111: M1r = 2'b01;
			14'b00100011100111: M1r = 2'b00;
			14'b01100011100111: M1r = 2'b01;
			14'b10100011100111: M1r = 2'b01;
			14'b11100011100111: M1r = 2'b01;
			14'b00110011100111: M1r = 2'b00;
			14'b01110011100111: M1r = 2'b00;
			14'b10110011100111: M1r = 2'b00;
			14'b11110011100111: M1r = 2'b00;
			14'b00000111100111: M1r = 2'b10;
			14'b01000111100111: M1r = 2'b10;
			14'b10000111100111: M1r = 2'b10;
			14'b11000111100111: M1r = 2'b11;
			14'b00010111100111: M1r = 2'b10;
			14'b01010111100111: M1r = 2'b10;
			14'b10010111100111: M1r = 2'b10;
			14'b11010111100111: M1r = 2'b10;
			14'b00100111100111: M1r = 2'b01;
			14'b01100111100111: M1r = 2'b01;
			14'b10100111100111: M1r = 2'b01;
			14'b11100111100111: M1r = 2'b10;
			14'b00110111100111: M1r = 2'b01;
			14'b01110111100111: M1r = 2'b01;
			14'b10110111100111: M1r = 2'b01;
			14'b11110111100111: M1r = 2'b01;
			14'b00001011100111: M1r = 2'b11;
			14'b01001011100111: M1r = 2'b11;
			14'b10001011100111: M1r = 2'b11;
			14'b11001011100111: M1r = 2'b11;
			14'b00011011100111: M1r = 2'b10;
			14'b01011011100111: M1r = 2'b10;
			14'b10011011100111: M1r = 2'b11;
			14'b11011011100111: M1r = 2'b11;
			14'b00101011100111: M1r = 2'b10;
			14'b01101011100111: M1r = 2'b10;
			14'b10101011100111: M1r = 2'b10;
			14'b11101011100111: M1r = 2'b10;
			14'b00111011100111: M1r = 2'b01;
			14'b01111011100111: M1r = 2'b10;
			14'b10111011100111: M1r = 2'b10;
			14'b11111011100111: M1r = 2'b10;
			14'b00001111100111: M1r = 2'b11;
			14'b01001111100111: M1r = 2'b11;
			14'b10001111100111: M1r = 2'b11;
			14'b11001111100111: M1r = 2'b11;
			14'b00011111100111: M1r = 2'b11;
			14'b01011111100111: M1r = 2'b11;
			14'b10011111100111: M1r = 2'b11;
			14'b11011111100111: M1r = 2'b11;
			14'b00101111100111: M1r = 2'b11;
			14'b01101111100111: M1r = 2'b11;
			14'b10101111100111: M1r = 2'b11;
			14'b11101111100111: M1r = 2'b11;
			14'b00111111100111: M1r = 2'b10;
			14'b01111111100111: M1r = 2'b10;
			14'b10111111100111: M1r = 2'b10;
			14'b11111111100111: M1r = 2'b11;
			14'b00000000110111: M1r = 2'b11;
			14'b01000000110111: M1r = 2'b11;
			14'b10000000110111: M1r = 2'b11;
			14'b11000000110111: M1r = 2'b11;
			14'b00010000110111: M1r = 2'b10;
			14'b01010000110111: M1r = 2'b10;
			14'b10010000110111: M1r = 2'b10;
			14'b11010000110111: M1r = 2'b11;
			14'b00100000110111: M1r = 2'b10;
			14'b01100000110111: M1r = 2'b10;
			14'b10100000110111: M1r = 2'b10;
			14'b11100000110111: M1r = 2'b10;
			14'b00110000110111: M1r = 2'b01;
			14'b01110000110111: M1r = 2'b01;
			14'b10110000110111: M1r = 2'b01;
			14'b11110000110111: M1r = 2'b10;
			14'b00000100110111: M1r = 2'b11;
			14'b01000100110111: M1r = 2'b11;
			14'b10000100110111: M1r = 2'b11;
			14'b11000100110111: M1r = 2'b11;
			14'b00010100110111: M1r = 2'b11;
			14'b01010100110111: M1r = 2'b11;
			14'b10010100110111: M1r = 2'b11;
			14'b11010100110111: M1r = 2'b11;
			14'b00100100110111: M1r = 2'b10;
			14'b01100100110111: M1r = 2'b11;
			14'b10100100110111: M1r = 2'b11;
			14'b11100100110111: M1r = 2'b11;
			14'b00110100110111: M1r = 2'b10;
			14'b01110100110111: M1r = 2'b10;
			14'b10110100110111: M1r = 2'b10;
			14'b11110100110111: M1r = 2'b10;
			14'b00001000110111: M1r = 2'b11;
			14'b01001000110111: M1r = 2'b11;
			14'b10001000110111: M1r = 2'b11;
			14'b11001000110111: M1r = 2'b11;
			14'b00011000110111: M1r = 2'b11;
			14'b01011000110111: M1r = 2'b11;
			14'b10011000110111: M1r = 2'b11;
			14'b11011000110111: M1r = 2'b11;
			14'b00101000110111: M1r = 2'b11;
			14'b01101000110111: M1r = 2'b11;
			14'b10101000110111: M1r = 2'b11;
			14'b11101000110111: M1r = 2'b11;
			14'b00111000110111: M1r = 2'b11;
			14'b01111000110111: M1r = 2'b11;
			14'b10111000110111: M1r = 2'b11;
			14'b11111000110111: M1r = 2'b11;
			14'b00001100110111: M1r = 2'b11;
			14'b01001100110111: M1r = 2'b11;
			14'b10001100110111: M1r = 2'b11;
			14'b11001100110111: M1r = 2'b11;
			14'b00011100110111: M1r = 2'b11;
			14'b01011100110111: M1r = 2'b11;
			14'b10011100110111: M1r = 2'b11;
			14'b11011100110111: M1r = 2'b11;
			14'b00101100110111: M1r = 2'b11;
			14'b01101100110111: M1r = 2'b11;
			14'b10101100110111: M1r = 2'b11;
			14'b11101100110111: M1r = 2'b11;
			14'b00111100110111: M1r = 2'b11;
			14'b01111100110111: M1r = 2'b11;
			14'b10111100110111: M1r = 2'b11;
			14'b11111100110111: M1r = 2'b11;
			14'b00000001110111: M1r = 2'b10;
			14'b01000001110111: M1r = 2'b10;
			14'b10000001110111: M1r = 2'b11;
			14'b11000001110111: M1r = 2'b11;
			14'b00010001110111: M1r = 2'b10;
			14'b01010001110111: M1r = 2'b10;
			14'b10010001110111: M1r = 2'b10;
			14'b11010001110111: M1r = 2'b10;
			14'b00100001110111: M1r = 2'b01;
			14'b01100001110111: M1r = 2'b01;
			14'b10100001110111: M1r = 2'b10;
			14'b11100001110111: M1r = 2'b10;
			14'b00110001110111: M1r = 2'b01;
			14'b01110001110111: M1r = 2'b01;
			14'b10110001110111: M1r = 2'b01;
			14'b11110001110111: M1r = 2'b01;
			14'b00000101110111: M1r = 2'b11;
			14'b01000101110111: M1r = 2'b11;
			14'b10000101110111: M1r = 2'b11;
			14'b11000101110111: M1r = 2'b11;
			14'b00010101110111: M1r = 2'b11;
			14'b01010101110111: M1r = 2'b11;
			14'b10010101110111: M1r = 2'b11;
			14'b11010101110111: M1r = 2'b11;
			14'b00100101110111: M1r = 2'b10;
			14'b01100101110111: M1r = 2'b10;
			14'b10100101110111: M1r = 2'b10;
			14'b11100101110111: M1r = 2'b11;
			14'b00110101110111: M1r = 2'b10;
			14'b01110101110111: M1r = 2'b10;
			14'b10110101110111: M1r = 2'b10;
			14'b11110101110111: M1r = 2'b10;
			14'b00001001110111: M1r = 2'b11;
			14'b01001001110111: M1r = 2'b11;
			14'b10001001110111: M1r = 2'b11;
			14'b11001001110111: M1r = 2'b11;
			14'b00011001110111: M1r = 2'b11;
			14'b01011001110111: M1r = 2'b11;
			14'b10011001110111: M1r = 2'b11;
			14'b11011001110111: M1r = 2'b11;
			14'b00101001110111: M1r = 2'b11;
			14'b01101001110111: M1r = 2'b11;
			14'b10101001110111: M1r = 2'b11;
			14'b11101001110111: M1r = 2'b11;
			14'b00111001110111: M1r = 2'b10;
			14'b01111001110111: M1r = 2'b11;
			14'b10111001110111: M1r = 2'b11;
			14'b11111001110111: M1r = 2'b11;
			14'b00001101110111: M1r = 2'b11;
			14'b01001101110111: M1r = 2'b11;
			14'b10001101110111: M1r = 2'b11;
			14'b11001101110111: M1r = 2'b11;
			14'b00011101110111: M1r = 2'b11;
			14'b01011101110111: M1r = 2'b11;
			14'b10011101110111: M1r = 2'b11;
			14'b11011101110111: M1r = 2'b11;
			14'b00101101110111: M1r = 2'b11;
			14'b01101101110111: M1r = 2'b11;
			14'b10101101110111: M1r = 2'b11;
			14'b11101101110111: M1r = 2'b11;
			14'b00111101110111: M1r = 2'b11;
			14'b01111101110111: M1r = 2'b11;
			14'b10111101110111: M1r = 2'b11;
			14'b11111101110111: M1r = 2'b11;
			14'b00000010110111: M1r = 2'b10;
			14'b01000010110111: M1r = 2'b10;
			14'b10000010110111: M1r = 2'b10;
			14'b11000010110111: M1r = 2'b10;
			14'b00010010110111: M1r = 2'b10;
			14'b01010010110111: M1r = 2'b10;
			14'b10010010110111: M1r = 2'b10;
			14'b11010010110111: M1r = 2'b10;
			14'b00100010110111: M1r = 2'b01;
			14'b01100010110111: M1r = 2'b01;
			14'b10100010110111: M1r = 2'b01;
			14'b11100010110111: M1r = 2'b10;
			14'b00110010110111: M1r = 2'b01;
			14'b01110010110111: M1r = 2'b01;
			14'b10110010110111: M1r = 2'b01;
			14'b11110010110111: M1r = 2'b01;
			14'b00000110110111: M1r = 2'b11;
			14'b01000110110111: M1r = 2'b11;
			14'b10000110110111: M1r = 2'b11;
			14'b11000110110111: M1r = 2'b11;
			14'b00010110110111: M1r = 2'b10;
			14'b01010110110111: M1r = 2'b10;
			14'b10010110110111: M1r = 2'b11;
			14'b11010110110111: M1r = 2'b11;
			14'b00100110110111: M1r = 2'b10;
			14'b01100110110111: M1r = 2'b10;
			14'b10100110110111: M1r = 2'b10;
			14'b11100110110111: M1r = 2'b10;
			14'b00110110110111: M1r = 2'b01;
			14'b01110110110111: M1r = 2'b01;
			14'b10110110110111: M1r = 2'b10;
			14'b11110110110111: M1r = 2'b10;
			14'b00001010110111: M1r = 2'b11;
			14'b01001010110111: M1r = 2'b11;
			14'b10001010110111: M1r = 2'b11;
			14'b11001010110111: M1r = 2'b11;
			14'b00011010110111: M1r = 2'b11;
			14'b01011010110111: M1r = 2'b11;
			14'b10011010110111: M1r = 2'b11;
			14'b11011010110111: M1r = 2'b11;
			14'b00101010110111: M1r = 2'b11;
			14'b01101010110111: M1r = 2'b11;
			14'b10101010110111: M1r = 2'b11;
			14'b11101010110111: M1r = 2'b11;
			14'b00111010110111: M1r = 2'b10;
			14'b01111010110111: M1r = 2'b10;
			14'b10111010110111: M1r = 2'b10;
			14'b11111010110111: M1r = 2'b11;
			14'b00001110110111: M1r = 2'b11;
			14'b01001110110111: M1r = 2'b11;
			14'b10001110110111: M1r = 2'b11;
			14'b11001110110111: M1r = 2'b11;
			14'b00011110110111: M1r = 2'b11;
			14'b01011110110111: M1r = 2'b11;
			14'b10011110110111: M1r = 2'b11;
			14'b11011110110111: M1r = 2'b11;
			14'b00101110110111: M1r = 2'b11;
			14'b01101110110111: M1r = 2'b11;
			14'b10101110110111: M1r = 2'b11;
			14'b11101110110111: M1r = 2'b11;
			14'b00111110110111: M1r = 2'b11;
			14'b01111110110111: M1r = 2'b11;
			14'b10111110110111: M1r = 2'b11;
			14'b11111110110111: M1r = 2'b11;
			14'b00000011110111: M1r = 2'b10;
			14'b01000011110111: M1r = 2'b10;
			14'b10000011110111: M1r = 2'b10;
			14'b11000011110111: M1r = 2'b10;
			14'b00010011110111: M1r = 2'b01;
			14'b01010011110111: M1r = 2'b01;
			14'b10010011110111: M1r = 2'b10;
			14'b11010011110111: M1r = 2'b10;
			14'b00100011110111: M1r = 2'b01;
			14'b01100011110111: M1r = 2'b01;
			14'b10100011110111: M1r = 2'b01;
			14'b11100011110111: M1r = 2'b01;
			14'b00110011110111: M1r = 2'b00;
			14'b01110011110111: M1r = 2'b00;
			14'b10110011110111: M1r = 2'b01;
			14'b11110011110111: M1r = 2'b01;
			14'b00000111110111: M1r = 2'b10;
			14'b01000111110111: M1r = 2'b11;
			14'b10000111110111: M1r = 2'b11;
			14'b11000111110111: M1r = 2'b11;
			14'b00010111110111: M1r = 2'b10;
			14'b01010111110111: M1r = 2'b10;
			14'b10010111110111: M1r = 2'b10;
			14'b11010111110111: M1r = 2'b10;
			14'b00100111110111: M1r = 2'b10;
			14'b01100111110111: M1r = 2'b10;
			14'b10100111110111: M1r = 2'b10;
			14'b11100111110111: M1r = 2'b10;
			14'b00110111110111: M1r = 2'b01;
			14'b01110111110111: M1r = 2'b01;
			14'b10110111110111: M1r = 2'b01;
			14'b11110111110111: M1r = 2'b10;
			14'b00001011110111: M1r = 2'b11;
			14'b01001011110111: M1r = 2'b11;
			14'b10001011110111: M1r = 2'b11;
			14'b11001011110111: M1r = 2'b11;
			14'b00011011110111: M1r = 2'b11;
			14'b01011011110111: M1r = 2'b11;
			14'b10011011110111: M1r = 2'b11;
			14'b11011011110111: M1r = 2'b11;
			14'b00101011110111: M1r = 2'b10;
			14'b01101011110111: M1r = 2'b10;
			14'b10101011110111: M1r = 2'b11;
			14'b11101011110111: M1r = 2'b11;
			14'b00111011110111: M1r = 2'b10;
			14'b01111011110111: M1r = 2'b10;
			14'b10111011110111: M1r = 2'b10;
			14'b11111011110111: M1r = 2'b10;
			14'b00001111110111: M1r = 2'b11;
			14'b01001111110111: M1r = 2'b11;
			14'b10001111110111: M1r = 2'b11;
			14'b11001111110111: M1r = 2'b11;
			14'b00011111110111: M1r = 2'b11;
			14'b01011111110111: M1r = 2'b11;
			14'b10011111110111: M1r = 2'b11;
			14'b11011111110111: M1r = 2'b11;
			14'b00101111110111: M1r = 2'b11;
			14'b01101111110111: M1r = 2'b11;
			14'b10101111110111: M1r = 2'b11;
			14'b11101111110111: M1r = 2'b11;
			14'b00111111110111: M1r = 2'b11;
			14'b01111111110111: M1r = 2'b11;
			14'b10111111110111: M1r = 2'b11;
			14'b11111111110111: M1r = 2'b11;
			14'b00000000001011: M1r = 2'b00;
			14'b01000000001011: M1r = 2'b01;
			14'b10000000001011: M1r = 2'b01;
			14'b11000000001011: M1r = 2'b01;
			14'b00010000001011: M1r = 2'b00;
			14'b01010000001011: M1r = 2'b00;
			14'b10010000001011: M1r = 2'b00;
			14'b11010000001011: M1r = 2'b00;
			14'b00100000001011: M1r = 2'b00;
			14'b01100000001011: M1r = 2'b00;
			14'b10100000001011: M1r = 2'b00;
			14'b11100000001011: M1r = 2'b00;
			14'b00110000001011: M1r = 2'b00;
			14'b01110000001011: M1r = 2'b00;
			14'b10110000001011: M1r = 2'b00;
			14'b11110000001011: M1r = 2'b00;
			14'b00000100001011: M1r = 2'b01;
			14'b01000100001011: M1r = 2'b01;
			14'b10000100001011: M1r = 2'b10;
			14'b11000100001011: M1r = 2'b10;
			14'b00010100001011: M1r = 2'b01;
			14'b01010100001011: M1r = 2'b01;
			14'b10010100001011: M1r = 2'b01;
			14'b11010100001011: M1r = 2'b01;
			14'b00100100001011: M1r = 2'b00;
			14'b01100100001011: M1r = 2'b00;
			14'b10100100001011: M1r = 2'b01;
			14'b11100100001011: M1r = 2'b01;
			14'b00110100001011: M1r = 2'b00;
			14'b01110100001011: M1r = 2'b00;
			14'b10110100001011: M1r = 2'b00;
			14'b11110100001011: M1r = 2'b00;
			14'b00001000001011: M1r = 2'b10;
			14'b01001000001011: M1r = 2'b10;
			14'b10001000001011: M1r = 2'b10;
			14'b11001000001011: M1r = 2'b10;
			14'b00011000001011: M1r = 2'b10;
			14'b01011000001011: M1r = 2'b10;
			14'b10011000001011: M1r = 2'b10;
			14'b11011000001011: M1r = 2'b10;
			14'b00101000001011: M1r = 2'b01;
			14'b01101000001011: M1r = 2'b01;
			14'b10101000001011: M1r = 2'b01;
			14'b11101000001011: M1r = 2'b10;
			14'b00111000001011: M1r = 2'b01;
			14'b01111000001011: M1r = 2'b01;
			14'b10111000001011: M1r = 2'b01;
			14'b11111000001011: M1r = 2'b01;
			14'b00001100001011: M1r = 2'b11;
			14'b01001100001011: M1r = 2'b11;
			14'b10001100001011: M1r = 2'b11;
			14'b11001100001011: M1r = 2'b11;
			14'b00011100001011: M1r = 2'b10;
			14'b01011100001011: M1r = 2'b10;
			14'b10011100001011: M1r = 2'b11;
			14'b11011100001011: M1r = 2'b11;
			14'b00101100001011: M1r = 2'b10;
			14'b01101100001011: M1r = 2'b10;
			14'b10101100001011: M1r = 2'b10;
			14'b11101100001011: M1r = 2'b10;
			14'b00111100001011: M1r = 2'b01;
			14'b01111100001011: M1r = 2'b01;
			14'b10111100001011: M1r = 2'b10;
			14'b11111100001011: M1r = 2'b10;
			14'b00000001001011: M1r = 2'b00;
			14'b01000001001011: M1r = 2'b00;
			14'b10000001001011: M1r = 2'b01;
			14'b11000001001011: M1r = 2'b01;
			14'b00010001001011: M1r = 2'b00;
			14'b01010001001011: M1r = 2'b00;
			14'b10010001001011: M1r = 2'b00;
			14'b11010001001011: M1r = 2'b00;
			14'b00100001001011: M1r = 2'b00;
			14'b01100001001011: M1r = 2'b00;
			14'b10100001001011: M1r = 2'b00;
			14'b11100001001011: M1r = 2'b00;
			14'b00110001001011: M1r = 2'b00;
			14'b01110001001011: M1r = 2'b00;
			14'b10110001001011: M1r = 2'b00;
			14'b11110001001011: M1r = 2'b00;
			14'b00000101001011: M1r = 2'b01;
			14'b01000101001011: M1r = 2'b01;
			14'b10000101001011: M1r = 2'b01;
			14'b11000101001011: M1r = 2'b01;
			14'b00010101001011: M1r = 2'b00;
			14'b01010101001011: M1r = 2'b01;
			14'b10010101001011: M1r = 2'b01;
			14'b11010101001011: M1r = 2'b01;
			14'b00100101001011: M1r = 2'b00;
			14'b01100101001011: M1r = 2'b00;
			14'b10100101001011: M1r = 2'b00;
			14'b11100101001011: M1r = 2'b00;
			14'b00110101001011: M1r = 2'b00;
			14'b01110101001011: M1r = 2'b00;
			14'b10110101001011: M1r = 2'b00;
			14'b11110101001011: M1r = 2'b00;
			14'b00001001001011: M1r = 2'b10;
			14'b01001001001011: M1r = 2'b10;
			14'b10001001001011: M1r = 2'b10;
			14'b11001001001011: M1r = 2'b10;
			14'b00011001001011: M1r = 2'b01;
			14'b01011001001011: M1r = 2'b01;
			14'b10011001001011: M1r = 2'b10;
			14'b11011001001011: M1r = 2'b10;
			14'b00101001001011: M1r = 2'b01;
			14'b01101001001011: M1r = 2'b01;
			14'b10101001001011: M1r = 2'b01;
			14'b11101001001011: M1r = 2'b01;
			14'b00111001001011: M1r = 2'b00;
			14'b01111001001011: M1r = 2'b00;
			14'b10111001001011: M1r = 2'b01;
			14'b11111001001011: M1r = 2'b01;
			14'b00001101001011: M1r = 2'b10;
			14'b01001101001011: M1r = 2'b11;
			14'b10001101001011: M1r = 2'b11;
			14'b11001101001011: M1r = 2'b11;
			14'b00011101001011: M1r = 2'b10;
			14'b01011101001011: M1r = 2'b10;
			14'b10011101001011: M1r = 2'b10;
			14'b11011101001011: M1r = 2'b10;
			14'b00101101001011: M1r = 2'b10;
			14'b01101101001011: M1r = 2'b10;
			14'b10101101001011: M1r = 2'b10;
			14'b11101101001011: M1r = 2'b10;
			14'b00111101001011: M1r = 2'b01;
			14'b01111101001011: M1r = 2'b01;
			14'b10111101001011: M1r = 2'b01;
			14'b11111101001011: M1r = 2'b10;
			14'b00000010001011: M1r = 2'b00;
			14'b01000010001011: M1r = 2'b00;
			14'b10000010001011: M1r = 2'b00;
			14'b11000010001011: M1r = 2'b00;
			14'b00010010001011: M1r = 2'b00;
			14'b01010010001011: M1r = 2'b00;
			14'b10010010001011: M1r = 2'b00;
			14'b11010010001011: M1r = 2'b00;
			14'b00100010001011: M1r = 2'b00;
			14'b01100010001011: M1r = 2'b00;
			14'b10100010001011: M1r = 2'b00;
			14'b11100010001011: M1r = 2'b00;
			14'b00110010001011: M1r = 2'b00;
			14'b01110010001011: M1r = 2'b00;
			14'b10110010001011: M1r = 2'b00;
			14'b11110010001011: M1r = 2'b00;
			14'b00000110001011: M1r = 2'b01;
			14'b01000110001011: M1r = 2'b01;
			14'b10000110001011: M1r = 2'b01;
			14'b11000110001011: M1r = 2'b01;
			14'b00010110001011: M1r = 2'b00;
			14'b01010110001011: M1r = 2'b00;
			14'b10010110001011: M1r = 2'b01;
			14'b11010110001011: M1r = 2'b01;
			14'b00100110001011: M1r = 2'b00;
			14'b01100110001011: M1r = 2'b00;
			14'b10100110001011: M1r = 2'b00;
			14'b11100110001011: M1r = 2'b00;
			14'b00110110001011: M1r = 2'b00;
			14'b01110110001011: M1r = 2'b00;
			14'b10110110001011: M1r = 2'b00;
			14'b11110110001011: M1r = 2'b00;
			14'b00001010001011: M1r = 2'b01;
			14'b01001010001011: M1r = 2'b10;
			14'b10001010001011: M1r = 2'b10;
			14'b11001010001011: M1r = 2'b10;
			14'b00011010001011: M1r = 2'b01;
			14'b01011010001011: M1r = 2'b01;
			14'b10011010001011: M1r = 2'b01;
			14'b11011010001011: M1r = 2'b01;
			14'b00101010001011: M1r = 2'b00;
			14'b01101010001011: M1r = 2'b01;
			14'b10101010001011: M1r = 2'b01;
			14'b11101010001011: M1r = 2'b01;
			14'b00111010001011: M1r = 2'b00;
			14'b01111010001011: M1r = 2'b00;
			14'b10111010001011: M1r = 2'b00;
			14'b11111010001011: M1r = 2'b00;
			14'b00001110001011: M1r = 2'b10;
			14'b01001110001011: M1r = 2'b10;
			14'b10001110001011: M1r = 2'b10;
			14'b11001110001011: M1r = 2'b11;
			14'b00011110001011: M1r = 2'b10;
			14'b01011110001011: M1r = 2'b10;
			14'b10011110001011: M1r = 2'b10;
			14'b11011110001011: M1r = 2'b10;
			14'b00101110001011: M1r = 2'b01;
			14'b01101110001011: M1r = 2'b01;
			14'b10101110001011: M1r = 2'b10;
			14'b11101110001011: M1r = 2'b10;
			14'b00111110001011: M1r = 2'b01;
			14'b01111110001011: M1r = 2'b01;
			14'b10111110001011: M1r = 2'b01;
			14'b11111110001011: M1r = 2'b01;
			14'b00000011001011: M1r = 2'b00;
			14'b01000011001011: M1r = 2'b00;
			14'b10000011001011: M1r = 2'b00;
			14'b11000011001011: M1r = 2'b00;
			14'b00010011001011: M1r = 2'b00;
			14'b01010011001011: M1r = 2'b00;
			14'b10010011001011: M1r = 2'b00;
			14'b11010011001011: M1r = 2'b00;
			14'b00100011001011: M1r = 2'b00;
			14'b01100011001011: M1r = 2'b00;
			14'b10100011001011: M1r = 2'b00;
			14'b11100011001011: M1r = 2'b00;
			14'b00110011001011: M1r = 2'b00;
			14'b01110011001011: M1r = 2'b00;
			14'b10110011001011: M1r = 2'b00;
			14'b11110011001011: M1r = 2'b00;
			14'b00000111001011: M1r = 2'b00;
			14'b01000111001011: M1r = 2'b01;
			14'b10000111001011: M1r = 2'b01;
			14'b11000111001011: M1r = 2'b01;
			14'b00010111001011: M1r = 2'b00;
			14'b01010111001011: M1r = 2'b00;
			14'b10010111001011: M1r = 2'b00;
			14'b11010111001011: M1r = 2'b00;
			14'b00100111001011: M1r = 2'b00;
			14'b01100111001011: M1r = 2'b00;
			14'b10100111001011: M1r = 2'b00;
			14'b11100111001011: M1r = 2'b00;
			14'b00110111001011: M1r = 2'b00;
			14'b01110111001011: M1r = 2'b00;
			14'b10110111001011: M1r = 2'b00;
			14'b11110111001011: M1r = 2'b00;
			14'b00001011001011: M1r = 2'b01;
			14'b01001011001011: M1r = 2'b01;
			14'b10001011001011: M1r = 2'b01;
			14'b11001011001011: M1r = 2'b10;
			14'b00011011001011: M1r = 2'b01;
			14'b01011011001011: M1r = 2'b01;
			14'b10011011001011: M1r = 2'b01;
			14'b11011011001011: M1r = 2'b01;
			14'b00101011001011: M1r = 2'b00;
			14'b01101011001011: M1r = 2'b00;
			14'b10101011001011: M1r = 2'b01;
			14'b11101011001011: M1r = 2'b01;
			14'b00111011001011: M1r = 2'b00;
			14'b01111011001011: M1r = 2'b00;
			14'b10111011001011: M1r = 2'b00;
			14'b11111011001011: M1r = 2'b00;
			14'b00001111001011: M1r = 2'b10;
			14'b01001111001011: M1r = 2'b10;
			14'b10001111001011: M1r = 2'b10;
			14'b11001111001011: M1r = 2'b10;
			14'b00011111001011: M1r = 2'b01;
			14'b01011111001011: M1r = 2'b10;
			14'b10011111001011: M1r = 2'b10;
			14'b11011111001011: M1r = 2'b10;
			14'b00101111001011: M1r = 2'b01;
			14'b01101111001011: M1r = 2'b01;
			14'b10101111001011: M1r = 2'b01;
			14'b11101111001011: M1r = 2'b01;
			14'b00111111001011: M1r = 2'b00;
			14'b01111111001011: M1r = 2'b01;
			14'b10111111001011: M1r = 2'b01;
			14'b11111111001011: M1r = 2'b01;
			14'b00000000011011: M1r = 2'b01;
			14'b01000000011011: M1r = 2'b01;
			14'b10000000011011: M1r = 2'b01;
			14'b11000000011011: M1r = 2'b01;
			14'b00010000011011: M1r = 2'b00;
			14'b01010000011011: M1r = 2'b01;
			14'b10010000011011: M1r = 2'b01;
			14'b11010000011011: M1r = 2'b01;
			14'b00100000011011: M1r = 2'b00;
			14'b01100000011011: M1r = 2'b00;
			14'b10100000011011: M1r = 2'b00;
			14'b11100000011011: M1r = 2'b00;
			14'b00110000011011: M1r = 2'b00;
			14'b01110000011011: M1r = 2'b00;
			14'b10110000011011: M1r = 2'b00;
			14'b11110000011011: M1r = 2'b00;
			14'b00000100011011: M1r = 2'b10;
			14'b01000100011011: M1r = 2'b10;
			14'b10000100011011: M1r = 2'b10;
			14'b11000100011011: M1r = 2'b10;
			14'b00010100011011: M1r = 2'b01;
			14'b01010100011011: M1r = 2'b01;
			14'b10010100011011: M1r = 2'b10;
			14'b11010100011011: M1r = 2'b10;
			14'b00100100011011: M1r = 2'b01;
			14'b01100100011011: M1r = 2'b01;
			14'b10100100011011: M1r = 2'b01;
			14'b11100100011011: M1r = 2'b01;
			14'b00110100011011: M1r = 2'b00;
			14'b01110100011011: M1r = 2'b00;
			14'b10110100011011: M1r = 2'b01;
			14'b11110100011011: M1r = 2'b01;
			14'b00001000011011: M1r = 2'b10;
			14'b01001000011011: M1r = 2'b11;
			14'b10001000011011: M1r = 2'b11;
			14'b11001000011011: M1r = 2'b11;
			14'b00011000011011: M1r = 2'b10;
			14'b01011000011011: M1r = 2'b10;
			14'b10011000011011: M1r = 2'b10;
			14'b11011000011011: M1r = 2'b10;
			14'b00101000011011: M1r = 2'b01;
			14'b01101000011011: M1r = 2'b10;
			14'b10101000011011: M1r = 2'b10;
			14'b11101000011011: M1r = 2'b10;
			14'b00111000011011: M1r = 2'b01;
			14'b01111000011011: M1r = 2'b01;
			14'b10111000011011: M1r = 2'b01;
			14'b11111000011011: M1r = 2'b01;
			14'b00001100011011: M1r = 2'b11;
			14'b01001100011011: M1r = 2'b11;
			14'b10001100011011: M1r = 2'b11;
			14'b11001100011011: M1r = 2'b11;
			14'b00011100011011: M1r = 2'b11;
			14'b01011100011011: M1r = 2'b11;
			14'b10011100011011: M1r = 2'b11;
			14'b11011100011011: M1r = 2'b11;
			14'b00101100011011: M1r = 2'b10;
			14'b01101100011011: M1r = 2'b10;
			14'b10101100011011: M1r = 2'b11;
			14'b11101100011011: M1r = 2'b11;
			14'b00111100011011: M1r = 2'b10;
			14'b01111100011011: M1r = 2'b10;
			14'b10111100011011: M1r = 2'b10;
			14'b11111100011011: M1r = 2'b10;
			14'b00000001011011: M1r = 2'b01;
			14'b01000001011011: M1r = 2'b01;
			14'b10000001011011: M1r = 2'b01;
			14'b11000001011011: M1r = 2'b01;
			14'b00010001011011: M1r = 2'b00;
			14'b01010001011011: M1r = 2'b00;
			14'b10010001011011: M1r = 2'b00;
			14'b11010001011011: M1r = 2'b01;
			14'b00100001011011: M1r = 2'b00;
			14'b01100001011011: M1r = 2'b00;
			14'b10100001011011: M1r = 2'b00;
			14'b11100001011011: M1r = 2'b00;
			14'b00110001011011: M1r = 2'b00;
			14'b01110001011011: M1r = 2'b00;
			14'b10110001011011: M1r = 2'b00;
			14'b11110001011011: M1r = 2'b00;
			14'b00000101011011: M1r = 2'b01;
			14'b01000101011011: M1r = 2'b10;
			14'b10000101011011: M1r = 2'b10;
			14'b11000101011011: M1r = 2'b10;
			14'b00010101011011: M1r = 2'b01;
			14'b01010101011011: M1r = 2'b01;
			14'b10010101011011: M1r = 2'b01;
			14'b11010101011011: M1r = 2'b01;
			14'b00100101011011: M1r = 2'b00;
			14'b01100101011011: M1r = 2'b01;
			14'b10100101011011: M1r = 2'b01;
			14'b11100101011011: M1r = 2'b01;
			14'b00110101011011: M1r = 2'b00;
			14'b01110101011011: M1r = 2'b00;
			14'b10110101011011: M1r = 2'b00;
			14'b11110101011011: M1r = 2'b00;
			14'b00001001011011: M1r = 2'b10;
			14'b01001001011011: M1r = 2'b10;
			14'b10001001011011: M1r = 2'b10;
			14'b11001001011011: M1r = 2'b11;
			14'b00011001011011: M1r = 2'b10;
			14'b01011001011011: M1r = 2'b10;
			14'b10011001011011: M1r = 2'b10;
			14'b11011001011011: M1r = 2'b10;
			14'b00101001011011: M1r = 2'b01;
			14'b01101001011011: M1r = 2'b01;
			14'b10101001011011: M1r = 2'b10;
			14'b11101001011011: M1r = 2'b10;
			14'b00111001011011: M1r = 2'b01;
			14'b01111001011011: M1r = 2'b01;
			14'b10111001011011: M1r = 2'b01;
			14'b11111001011011: M1r = 2'b01;
			14'b00001101011011: M1r = 2'b11;
			14'b01001101011011: M1r = 2'b11;
			14'b10001101011011: M1r = 2'b11;
			14'b11001101011011: M1r = 2'b11;
			14'b00011101011011: M1r = 2'b10;
			14'b01011101011011: M1r = 2'b11;
			14'b10011101011011: M1r = 2'b11;
			14'b11011101011011: M1r = 2'b11;
			14'b00101101011011: M1r = 2'b10;
			14'b01101101011011: M1r = 2'b10;
			14'b10101101011011: M1r = 2'b10;
			14'b11101101011011: M1r = 2'b10;
			14'b00111101011011: M1r = 2'b01;
			14'b01111101011011: M1r = 2'b10;
			14'b10111101011011: M1r = 2'b10;
			14'b11111101011011: M1r = 2'b10;
			14'b00000010011011: M1r = 2'b00;
			14'b01000010011011: M1r = 2'b01;
			14'b10000010011011: M1r = 2'b01;
			14'b11000010011011: M1r = 2'b01;
			14'b00010010011011: M1r = 2'b00;
			14'b01010010011011: M1r = 2'b00;
			14'b10010010011011: M1r = 2'b00;
			14'b11010010011011: M1r = 2'b00;
			14'b00100010011011: M1r = 2'b00;
			14'b01100010011011: M1r = 2'b00;
			14'b10100010011011: M1r = 2'b00;
			14'b11100010011011: M1r = 2'b00;
			14'b00110010011011: M1r = 2'b00;
			14'b01110010011011: M1r = 2'b00;
			14'b10110010011011: M1r = 2'b00;
			14'b11110010011011: M1r = 2'b00;
			14'b00000110011011: M1r = 2'b01;
			14'b01000110011011: M1r = 2'b01;
			14'b10000110011011: M1r = 2'b01;
			14'b11000110011011: M1r = 2'b10;
			14'b00010110011011: M1r = 2'b01;
			14'b01010110011011: M1r = 2'b01;
			14'b10010110011011: M1r = 2'b01;
			14'b11010110011011: M1r = 2'b01;
			14'b00100110011011: M1r = 2'b00;
			14'b01100110011011: M1r = 2'b00;
			14'b10100110011011: M1r = 2'b00;
			14'b11100110011011: M1r = 2'b01;
			14'b00110110011011: M1r = 2'b00;
			14'b01110110011011: M1r = 2'b00;
			14'b10110110011011: M1r = 2'b00;
			14'b11110110011011: M1r = 2'b00;
			14'b00001010011011: M1r = 2'b10;
			14'b01001010011011: M1r = 2'b10;
			14'b10001010011011: M1r = 2'b10;
			14'b11001010011011: M1r = 2'b10;
			14'b00011010011011: M1r = 2'b01;
			14'b01011010011011: M1r = 2'b10;
			14'b10011010011011: M1r = 2'b10;
			14'b11011010011011: M1r = 2'b10;
			14'b00101010011011: M1r = 2'b01;
			14'b01101010011011: M1r = 2'b01;
			14'b10101010011011: M1r = 2'b01;
			14'b11101010011011: M1r = 2'b01;
			14'b00111010011011: M1r = 2'b00;
			14'b01111010011011: M1r = 2'b01;
			14'b10111010011011: M1r = 2'b01;
			14'b11111010011011: M1r = 2'b01;
			14'b00001110011011: M1r = 2'b11;
			14'b01001110011011: M1r = 2'b11;
			14'b10001110011011: M1r = 2'b11;
			14'b11001110011011: M1r = 2'b11;
			14'b00011110011011: M1r = 2'b10;
			14'b01011110011011: M1r = 2'b10;
			14'b10011110011011: M1r = 2'b10;
			14'b11011110011011: M1r = 2'b11;
			14'b00101110011011: M1r = 2'b10;
			14'b01101110011011: M1r = 2'b10;
			14'b10101110011011: M1r = 2'b10;
			14'b11101110011011: M1r = 2'b10;
			14'b00111110011011: M1r = 2'b01;
			14'b01111110011011: M1r = 2'b01;
			14'b10111110011011: M1r = 2'b10;
			14'b11111110011011: M1r = 2'b10;
			14'b00000011011011: M1r = 2'b00;
			14'b01000011011011: M1r = 2'b00;
			14'b10000011011011: M1r = 2'b00;
			14'b11000011011011: M1r = 2'b01;
			14'b00010011011011: M1r = 2'b00;
			14'b01010011011011: M1r = 2'b00;
			14'b10010011011011: M1r = 2'b00;
			14'b11010011011011: M1r = 2'b00;
			14'b00100011011011: M1r = 2'b00;
			14'b01100011011011: M1r = 2'b00;
			14'b10100011011011: M1r = 2'b00;
			14'b11100011011011: M1r = 2'b00;
			14'b00110011011011: M1r = 2'b00;
			14'b01110011011011: M1r = 2'b00;
			14'b10110011011011: M1r = 2'b00;
			14'b11110011011011: M1r = 2'b00;
			14'b00000111011011: M1r = 2'b01;
			14'b01000111011011: M1r = 2'b01;
			14'b10000111011011: M1r = 2'b01;
			14'b11000111011011: M1r = 2'b01;
			14'b00010111011011: M1r = 2'b00;
			14'b01010111011011: M1r = 2'b01;
			14'b10010111011011: M1r = 2'b01;
			14'b11010111011011: M1r = 2'b01;
			14'b00100111011011: M1r = 2'b00;
			14'b01100111011011: M1r = 2'b00;
			14'b10100111011011: M1r = 2'b00;
			14'b11100111011011: M1r = 2'b00;
			14'b00110111011011: M1r = 2'b00;
			14'b01110111011011: M1r = 2'b00;
			14'b10110111011011: M1r = 2'b00;
			14'b11110111011011: M1r = 2'b00;
			14'b00001011011011: M1r = 2'b10;
			14'b01001011011011: M1r = 2'b10;
			14'b10001011011011: M1r = 2'b10;
			14'b11001011011011: M1r = 2'b10;
			14'b00011011011011: M1r = 2'b01;
			14'b01011011011011: M1r = 2'b01;
			14'b10011011011011: M1r = 2'b01;
			14'b11011011011011: M1r = 2'b10;
			14'b00101011011011: M1r = 2'b01;
			14'b01101011011011: M1r = 2'b01;
			14'b10101011011011: M1r = 2'b01;
			14'b11101011011011: M1r = 2'b01;
			14'b00111011011011: M1r = 2'b00;
			14'b01111011011011: M1r = 2'b00;
			14'b10111011011011: M1r = 2'b00;
			14'b11111011011011: M1r = 2'b01;
			14'b00001111011011: M1r = 2'b10;
			14'b01001111011011: M1r = 2'b10;
			14'b10001111011011: M1r = 2'b11;
			14'b11001111011011: M1r = 2'b11;
			14'b00011111011011: M1r = 2'b10;
			14'b01011111011011: M1r = 2'b10;
			14'b10011111011011: M1r = 2'b10;
			14'b11011111011011: M1r = 2'b10;
			14'b00101111011011: M1r = 2'b01;
			14'b01101111011011: M1r = 2'b10;
			14'b10101111011011: M1r = 2'b10;
			14'b11101111011011: M1r = 2'b10;
			14'b00111111011011: M1r = 2'b01;
			14'b01111111011011: M1r = 2'b01;
			14'b10111111011011: M1r = 2'b01;
			14'b11111111011011: M1r = 2'b01;
			14'b00000000101011: M1r = 2'b01;
			14'b01000000101011: M1r = 2'b10;
			14'b10000000101011: M1r = 2'b10;
			14'b11000000101011: M1r = 2'b10;
			14'b00010000101011: M1r = 2'b01;
			14'b01010000101011: M1r = 2'b01;
			14'b10010000101011: M1r = 2'b01;
			14'b11010000101011: M1r = 2'b01;
			14'b00100000101011: M1r = 2'b00;
			14'b01100000101011: M1r = 2'b01;
			14'b10100000101011: M1r = 2'b01;
			14'b11100000101011: M1r = 2'b01;
			14'b00110000101011: M1r = 2'b00;
			14'b01110000101011: M1r = 2'b00;
			14'b10110000101011: M1r = 2'b00;
			14'b11110000101011: M1r = 2'b00;
			14'b00000100101011: M1r = 2'b10;
			14'b01000100101011: M1r = 2'b10;
			14'b10000100101011: M1r = 2'b10;
			14'b11000100101011: M1r = 2'b11;
			14'b00010100101011: M1r = 2'b10;
			14'b01010100101011: M1r = 2'b10;
			14'b10010100101011: M1r = 2'b10;
			14'b11010100101011: M1r = 2'b10;
			14'b00100100101011: M1r = 2'b01;
			14'b01100100101011: M1r = 2'b01;
			14'b10100100101011: M1r = 2'b01;
			14'b11100100101011: M1r = 2'b10;
			14'b00110100101011: M1r = 2'b01;
			14'b01110100101011: M1r = 2'b01;
			14'b10110100101011: M1r = 2'b01;
			14'b11110100101011: M1r = 2'b01;
			14'b00001000101011: M1r = 2'b11;
			14'b01001000101011: M1r = 2'b11;
			14'b10001000101011: M1r = 2'b11;
			14'b11001000101011: M1r = 2'b11;
			14'b00011000101011: M1r = 2'b10;
			14'b01011000101011: M1r = 2'b11;
			14'b10011000101011: M1r = 2'b11;
			14'b11011000101011: M1r = 2'b11;
			14'b00101000101011: M1r = 2'b10;
			14'b01101000101011: M1r = 2'b10;
			14'b10101000101011: M1r = 2'b10;
			14'b11101000101011: M1r = 2'b10;
			14'b00111000101011: M1r = 2'b01;
			14'b01111000101011: M1r = 2'b10;
			14'b10111000101011: M1r = 2'b10;
			14'b11111000101011: M1r = 2'b10;
			14'b00001100101011: M1r = 2'b11;
			14'b01001100101011: M1r = 2'b11;
			14'b10001100101011: M1r = 2'b11;
			14'b11001100101011: M1r = 2'b11;
			14'b00011100101011: M1r = 2'b11;
			14'b01011100101011: M1r = 2'b11;
			14'b10011100101011: M1r = 2'b11;
			14'b11011100101011: M1r = 2'b11;
			14'b00101100101011: M1r = 2'b11;
			14'b01101100101011: M1r = 2'b11;
			14'b10101100101011: M1r = 2'b11;
			14'b11101100101011: M1r = 2'b11;
			14'b00111100101011: M1r = 2'b10;
			14'b01111100101011: M1r = 2'b10;
			14'b10111100101011: M1r = 2'b10;
			14'b11111100101011: M1r = 2'b11;
			14'b00000001101011: M1r = 2'b01;
			14'b01000001101011: M1r = 2'b01;
			14'b10000001101011: M1r = 2'b01;
			14'b11000001101011: M1r = 2'b10;
			14'b00010001101011: M1r = 2'b01;
			14'b01010001101011: M1r = 2'b01;
			14'b10010001101011: M1r = 2'b01;
			14'b11010001101011: M1r = 2'b01;
			14'b00100001101011: M1r = 2'b00;
			14'b01100001101011: M1r = 2'b00;
			14'b10100001101011: M1r = 2'b00;
			14'b11100001101011: M1r = 2'b01;
			14'b00110001101011: M1r = 2'b00;
			14'b01110001101011: M1r = 2'b00;
			14'b10110001101011: M1r = 2'b00;
			14'b11110001101011: M1r = 2'b00;
			14'b00000101101011: M1r = 2'b10;
			14'b01000101101011: M1r = 2'b10;
			14'b10000101101011: M1r = 2'b10;
			14'b11000101101011: M1r = 2'b10;
			14'b00010101101011: M1r = 2'b01;
			14'b01010101101011: M1r = 2'b10;
			14'b10010101101011: M1r = 2'b10;
			14'b11010101101011: M1r = 2'b10;
			14'b00100101101011: M1r = 2'b01;
			14'b01100101101011: M1r = 2'b01;
			14'b10100101101011: M1r = 2'b01;
			14'b11100101101011: M1r = 2'b01;
			14'b00110101101011: M1r = 2'b00;
			14'b01110101101011: M1r = 2'b01;
			14'b10110101101011: M1r = 2'b01;
			14'b11110101101011: M1r = 2'b01;
			14'b00001001101011: M1r = 2'b11;
			14'b01001001101011: M1r = 2'b11;
			14'b10001001101011: M1r = 2'b11;
			14'b11001001101011: M1r = 2'b11;
			14'b00011001101011: M1r = 2'b10;
			14'b01011001101011: M1r = 2'b10;
			14'b10011001101011: M1r = 2'b10;
			14'b11011001101011: M1r = 2'b11;
			14'b00101001101011: M1r = 2'b10;
			14'b01101001101011: M1r = 2'b10;
			14'b10101001101011: M1r = 2'b10;
			14'b11101001101011: M1r = 2'b10;
			14'b00111001101011: M1r = 2'b01;
			14'b01111001101011: M1r = 2'b01;
			14'b10111001101011: M1r = 2'b01;
			14'b11111001101011: M1r = 2'b10;
			14'b00001101101011: M1r = 2'b11;
			14'b01001101101011: M1r = 2'b11;
			14'b10001101101011: M1r = 2'b11;
			14'b11001101101011: M1r = 2'b11;
			14'b00011101101011: M1r = 2'b11;
			14'b01011101101011: M1r = 2'b11;
			14'b10011101101011: M1r = 2'b11;
			14'b11011101101011: M1r = 2'b11;
			14'b00101101101011: M1r = 2'b10;
			14'b01101101101011: M1r = 2'b11;
			14'b10101101101011: M1r = 2'b11;
			14'b11101101101011: M1r = 2'b11;
			14'b00111101101011: M1r = 2'b10;
			14'b01111101101011: M1r = 2'b10;
			14'b10111101101011: M1r = 2'b10;
			14'b11111101101011: M1r = 2'b10;
			14'b00000010101011: M1r = 2'b01;
			14'b01000010101011: M1r = 2'b01;
			14'b10000010101011: M1r = 2'b01;
			14'b11000010101011: M1r = 2'b01;
			14'b00010010101011: M1r = 2'b00;
			14'b01010010101011: M1r = 2'b00;
			14'b10010010101011: M1r = 2'b01;
			14'b11010010101011: M1r = 2'b01;
			14'b00100010101011: M1r = 2'b00;
			14'b01100010101011: M1r = 2'b00;
			14'b10100010101011: M1r = 2'b00;
			14'b11100010101011: M1r = 2'b00;
			14'b00110010101011: M1r = 2'b00;
			14'b01110010101011: M1r = 2'b00;
			14'b10110010101011: M1r = 2'b00;
			14'b11110010101011: M1r = 2'b00;
			14'b00000110101011: M1r = 2'b10;
			14'b01000110101011: M1r = 2'b10;
			14'b10000110101011: M1r = 2'b10;
			14'b11000110101011: M1r = 2'b10;
			14'b00010110101011: M1r = 2'b01;
			14'b01010110101011: M1r = 2'b01;
			14'b10010110101011: M1r = 2'b01;
			14'b11010110101011: M1r = 2'b10;
			14'b00100110101011: M1r = 2'b01;
			14'b01100110101011: M1r = 2'b01;
			14'b10100110101011: M1r = 2'b01;
			14'b11100110101011: M1r = 2'b01;
			14'b00110110101011: M1r = 2'b00;
			14'b01110110101011: M1r = 2'b00;
			14'b10110110101011: M1r = 2'b00;
			14'b11110110101011: M1r = 2'b01;
			14'b00001010101011: M1r = 2'b10;
			14'b01001010101011: M1r = 2'b10;
			14'b10001010101011: M1r = 2'b11;
			14'b11001010101011: M1r = 2'b11;
			14'b00011010101011: M1r = 2'b10;
			14'b01011010101011: M1r = 2'b10;
			14'b10011010101011: M1r = 2'b10;
			14'b11011010101011: M1r = 2'b10;
			14'b00101010101011: M1r = 2'b01;
			14'b01101010101011: M1r = 2'b10;
			14'b10101010101011: M1r = 2'b10;
			14'b11101010101011: M1r = 2'b10;
			14'b00111010101011: M1r = 2'b01;
			14'b01111010101011: M1r = 2'b01;
			14'b10111010101011: M1r = 2'b01;
			14'b11111010101011: M1r = 2'b01;
			14'b00001110101011: M1r = 2'b11;
			14'b01001110101011: M1r = 2'b11;
			14'b10001110101011: M1r = 2'b11;
			14'b11001110101011: M1r = 2'b11;
			14'b00011110101011: M1r = 2'b11;
			14'b01011110101011: M1r = 2'b11;
			14'b10011110101011: M1r = 2'b11;
			14'b11011110101011: M1r = 2'b11;
			14'b00101110101011: M1r = 2'b10;
			14'b01101110101011: M1r = 2'b10;
			14'b10101110101011: M1r = 2'b10;
			14'b11101110101011: M1r = 2'b11;
			14'b00111110101011: M1r = 2'b10;
			14'b01111110101011: M1r = 2'b10;
			14'b10111110101011: M1r = 2'b10;
			14'b11111110101011: M1r = 2'b10;
			14'b00000011101011: M1r = 2'b01;
			14'b01000011101011: M1r = 2'b01;
			14'b10000011101011: M1r = 2'b01;
			14'b11000011101011: M1r = 2'b01;
			14'b00010011101011: M1r = 2'b00;
			14'b01010011101011: M1r = 2'b00;
			14'b10010011101011: M1r = 2'b00;
			14'b11010011101011: M1r = 2'b01;
			14'b00100011101011: M1r = 2'b00;
			14'b01100011101011: M1r = 2'b00;
			14'b10100011101011: M1r = 2'b00;
			14'b11100011101011: M1r = 2'b00;
			14'b00110011101011: M1r = 2'b00;
			14'b01110011101011: M1r = 2'b00;
			14'b10110011101011: M1r = 2'b00;
			14'b11110011101011: M1r = 2'b00;
			14'b00000111101011: M1r = 2'b01;
			14'b01000111101011: M1r = 2'b01;
			14'b10000111101011: M1r = 2'b10;
			14'b11000111101011: M1r = 2'b10;
			14'b00010111101011: M1r = 2'b01;
			14'b01010111101011: M1r = 2'b01;
			14'b10010111101011: M1r = 2'b01;
			14'b11010111101011: M1r = 2'b01;
			14'b00100111101011: M1r = 2'b00;
			14'b01100111101011: M1r = 2'b00;
			14'b10100111101011: M1r = 2'b01;
			14'b11100111101011: M1r = 2'b01;
			14'b00110111101011: M1r = 2'b00;
			14'b01110111101011: M1r = 2'b00;
			14'b10110111101011: M1r = 2'b00;
			14'b11110111101011: M1r = 2'b00;
			14'b00001011101011: M1r = 2'b10;
			14'b01001011101011: M1r = 2'b10;
			14'b10001011101011: M1r = 2'b10;
			14'b11001011101011: M1r = 2'b10;
			14'b00011011101011: M1r = 2'b10;
			14'b01011011101011: M1r = 2'b10;
			14'b10011011101011: M1r = 2'b10;
			14'b11011011101011: M1r = 2'b10;
			14'b00101011101011: M1r = 2'b01;
			14'b01101011101011: M1r = 2'b01;
			14'b10101011101011: M1r = 2'b01;
			14'b11101011101011: M1r = 2'b10;
			14'b00111011101011: M1r = 2'b01;
			14'b01111011101011: M1r = 2'b01;
			14'b10111011101011: M1r = 2'b01;
			14'b11111011101011: M1r = 2'b01;
			14'b00001111101011: M1r = 2'b11;
			14'b01001111101011: M1r = 2'b11;
			14'b10001111101011: M1r = 2'b11;
			14'b11001111101011: M1r = 2'b11;
			14'b00011111101011: M1r = 2'b10;
			14'b01011111101011: M1r = 2'b10;
			14'b10011111101011: M1r = 2'b11;
			14'b11011111101011: M1r = 2'b11;
			14'b00101111101011: M1r = 2'b10;
			14'b01101111101011: M1r = 2'b10;
			14'b10101111101011: M1r = 2'b10;
			14'b11101111101011: M1r = 2'b10;
			14'b00111111101011: M1r = 2'b01;
			14'b01111111101011: M1r = 2'b10;
			14'b10111111101011: M1r = 2'b10;
			14'b11111111101011: M1r = 2'b10;
			14'b00000000111011: M1r = 2'b10;
			14'b01000000111011: M1r = 2'b10;
			14'b10000000111011: M1r = 2'b10;
			14'b11000000111011: M1r = 2'b10;
			14'b00010000111011: M1r = 2'b01;
			14'b01010000111011: M1r = 2'b01;
			14'b10010000111011: M1r = 2'b10;
			14'b11010000111011: M1r = 2'b10;
			14'b00100000111011: M1r = 2'b01;
			14'b01100000111011: M1r = 2'b01;
			14'b10100000111011: M1r = 2'b01;
			14'b11100000111011: M1r = 2'b01;
			14'b00110000111011: M1r = 2'b00;
			14'b01110000111011: M1r = 2'b01;
			14'b10110000111011: M1r = 2'b01;
			14'b11110000111011: M1r = 2'b01;
			14'b00000100111011: M1r = 2'b11;
			14'b01000100111011: M1r = 2'b11;
			14'b10000100111011: M1r = 2'b11;
			14'b11000100111011: M1r = 2'b11;
			14'b00010100111011: M1r = 2'b10;
			14'b01010100111011: M1r = 2'b10;
			14'b10010100111011: M1r = 2'b10;
			14'b11010100111011: M1r = 2'b11;
			14'b00100100111011: M1r = 2'b10;
			14'b01100100111011: M1r = 2'b10;
			14'b10100100111011: M1r = 2'b10;
			14'b11100100111011: M1r = 2'b10;
			14'b00110100111011: M1r = 2'b01;
			14'b01110100111011: M1r = 2'b01;
			14'b10110100111011: M1r = 2'b01;
			14'b11110100111011: M1r = 2'b10;
			14'b00001000111011: M1r = 2'b11;
			14'b01001000111011: M1r = 2'b11;
			14'b10001000111011: M1r = 2'b11;
			14'b11001000111011: M1r = 2'b11;
			14'b00011000111011: M1r = 2'b11;
			14'b01011000111011: M1r = 2'b11;
			14'b10011000111011: M1r = 2'b11;
			14'b11011000111011: M1r = 2'b11;
			14'b00101000111011: M1r = 2'b10;
			14'b01101000111011: M1r = 2'b10;
			14'b10101000111011: M1r = 2'b11;
			14'b11101000111011: M1r = 2'b11;
			14'b00111000111011: M1r = 2'b10;
			14'b01111000111011: M1r = 2'b10;
			14'b10111000111011: M1r = 2'b10;
			14'b11111000111011: M1r = 2'b10;
			14'b00001100111011: M1r = 2'b11;
			14'b01001100111011: M1r = 2'b11;
			14'b10001100111011: M1r = 2'b11;
			14'b11001100111011: M1r = 2'b11;
			14'b00011100111011: M1r = 2'b11;
			14'b01011100111011: M1r = 2'b11;
			14'b10011100111011: M1r = 2'b11;
			14'b11011100111011: M1r = 2'b11;
			14'b00101100111011: M1r = 2'b11;
			14'b01101100111011: M1r = 2'b11;
			14'b10101100111011: M1r = 2'b11;
			14'b11101100111011: M1r = 2'b11;
			14'b00111100111011: M1r = 2'b11;
			14'b01111100111011: M1r = 2'b11;
			14'b10111100111011: M1r = 2'b11;
			14'b11111100111011: M1r = 2'b11;
			14'b00000001111011: M1r = 2'b10;
			14'b01000001111011: M1r = 2'b10;
			14'b10000001111011: M1r = 2'b10;
			14'b11000001111011: M1r = 2'b10;
			14'b00010001111011: M1r = 2'b01;
			14'b01010001111011: M1r = 2'b01;
			14'b10010001111011: M1r = 2'b01;
			14'b11010001111011: M1r = 2'b01;
			14'b00100001111011: M1r = 2'b01;
			14'b01100001111011: M1r = 2'b01;
			14'b10100001111011: M1r = 2'b01;
			14'b11100001111011: M1r = 2'b01;
			14'b00110001111011: M1r = 2'b00;
			14'b01110001111011: M1r = 2'b00;
			14'b10110001111011: M1r = 2'b00;
			14'b11110001111011: M1r = 2'b01;
			14'b00000101111011: M1r = 2'b10;
			14'b01000101111011: M1r = 2'b10;
			14'b10000101111011: M1r = 2'b11;
			14'b11000101111011: M1r = 2'b11;
			14'b00010101111011: M1r = 2'b10;
			14'b01010101111011: M1r = 2'b10;
			14'b10010101111011: M1r = 2'b10;
			14'b11010101111011: M1r = 2'b10;
			14'b00100101111011: M1r = 2'b01;
			14'b01100101111011: M1r = 2'b01;
			14'b10100101111011: M1r = 2'b10;
			14'b11100101111011: M1r = 2'b10;
			14'b00110101111011: M1r = 2'b01;
			14'b01110101111011: M1r = 2'b01;
			14'b10110101111011: M1r = 2'b01;
			14'b11110101111011: M1r = 2'b01;
			14'b00001001111011: M1r = 2'b11;
			14'b01001001111011: M1r = 2'b11;
			14'b10001001111011: M1r = 2'b11;
			14'b11001001111011: M1r = 2'b11;
			14'b00011001111011: M1r = 2'b11;
			14'b01011001111011: M1r = 2'b11;
			14'b10011001111011: M1r = 2'b11;
			14'b11011001111011: M1r = 2'b11;
			14'b00101001111011: M1r = 2'b10;
			14'b01101001111011: M1r = 2'b10;
			14'b10101001111011: M1r = 2'b10;
			14'b11101001111011: M1r = 2'b11;
			14'b00111001111011: M1r = 2'b10;
			14'b01111001111011: M1r = 2'b10;
			14'b10111001111011: M1r = 2'b10;
			14'b11111001111011: M1r = 2'b10;
			14'b00001101111011: M1r = 2'b11;
			14'b01001101111011: M1r = 2'b11;
			14'b10001101111011: M1r = 2'b11;
			14'b11001101111011: M1r = 2'b11;
			14'b00011101111011: M1r = 2'b11;
			14'b01011101111011: M1r = 2'b11;
			14'b10011101111011: M1r = 2'b11;
			14'b11011101111011: M1r = 2'b11;
			14'b00101101111011: M1r = 2'b11;
			14'b01101101111011: M1r = 2'b11;
			14'b10101101111011: M1r = 2'b11;
			14'b11101101111011: M1r = 2'b11;
			14'b00111101111011: M1r = 2'b10;
			14'b01111101111011: M1r = 2'b10;
			14'b10111101111011: M1r = 2'b11;
			14'b11111101111011: M1r = 2'b11;
			14'b00000010111011: M1r = 2'b01;
			14'b01000010111011: M1r = 2'b01;
			14'b10000010111011: M1r = 2'b10;
			14'b11000010111011: M1r = 2'b10;
			14'b00010010111011: M1r = 2'b01;
			14'b01010010111011: M1r = 2'b01;
			14'b10010010111011: M1r = 2'b01;
			14'b11010010111011: M1r = 2'b01;
			14'b00100010111011: M1r = 2'b00;
			14'b01100010111011: M1r = 2'b00;
			14'b10100010111011: M1r = 2'b01;
			14'b11100010111011: M1r = 2'b01;
			14'b00110010111011: M1r = 2'b00;
			14'b01110010111011: M1r = 2'b00;
			14'b10110010111011: M1r = 2'b00;
			14'b11110010111011: M1r = 2'b00;
			14'b00000110111011: M1r = 2'b10;
			14'b01000110111011: M1r = 2'b10;
			14'b10000110111011: M1r = 2'b10;
			14'b11000110111011: M1r = 2'b10;
			14'b00010110111011: M1r = 2'b10;
			14'b01010110111011: M1r = 2'b10;
			14'b10010110111011: M1r = 2'b10;
			14'b11010110111011: M1r = 2'b10;
			14'b00100110111011: M1r = 2'b01;
			14'b01100110111011: M1r = 2'b01;
			14'b10100110111011: M1r = 2'b01;
			14'b11100110111011: M1r = 2'b01;
			14'b00110110111011: M1r = 2'b01;
			14'b01110110111011: M1r = 2'b01;
			14'b10110110111011: M1r = 2'b01;
			14'b11110110111011: M1r = 2'b01;
			14'b00001010111011: M1r = 2'b11;
			14'b01001010111011: M1r = 2'b11;
			14'b10001010111011: M1r = 2'b11;
			14'b11001010111011: M1r = 2'b11;
			14'b00011010111011: M1r = 2'b10;
			14'b01011010111011: M1r = 2'b10;
			14'b10011010111011: M1r = 2'b11;
			14'b11011010111011: M1r = 2'b11;
			14'b00101010111011: M1r = 2'b10;
			14'b01101010111011: M1r = 2'b10;
			14'b10101010111011: M1r = 2'b10;
			14'b11101010111011: M1r = 2'b10;
			14'b00111010111011: M1r = 2'b01;
			14'b01111010111011: M1r = 2'b01;
			14'b10111010111011: M1r = 2'b10;
			14'b11111010111011: M1r = 2'b10;
			14'b00001110111011: M1r = 2'b11;
			14'b01001110111011: M1r = 2'b11;
			14'b10001110111011: M1r = 2'b11;
			14'b11001110111011: M1r = 2'b11;
			14'b00011110111011: M1r = 2'b11;
			14'b01011110111011: M1r = 2'b11;
			14'b10011110111011: M1r = 2'b11;
			14'b11011110111011: M1r = 2'b11;
			14'b00101110111011: M1r = 2'b11;
			14'b01101110111011: M1r = 2'b11;
			14'b10101110111011: M1r = 2'b11;
			14'b11101110111011: M1r = 2'b11;
			14'b00111110111011: M1r = 2'b10;
			14'b01111110111011: M1r = 2'b10;
			14'b10111110111011: M1r = 2'b10;
			14'b11111110111011: M1r = 2'b11;
			14'b00000011111011: M1r = 2'b01;
			14'b01000011111011: M1r = 2'b01;
			14'b10000011111011: M1r = 2'b01;
			14'b11000011111011: M1r = 2'b01;
			14'b00010011111011: M1r = 2'b00;
			14'b01010011111011: M1r = 2'b01;
			14'b10010011111011: M1r = 2'b01;
			14'b11010011111011: M1r = 2'b01;
			14'b00100011111011: M1r = 2'b00;
			14'b01100011111011: M1r = 2'b00;
			14'b10100011111011: M1r = 2'b00;
			14'b11100011111011: M1r = 2'b00;
			14'b00110011111011: M1r = 2'b00;
			14'b01110011111011: M1r = 2'b00;
			14'b10110011111011: M1r = 2'b00;
			14'b11110011111011: M1r = 2'b00;
			14'b00000111111011: M1r = 2'b10;
			14'b01000111111011: M1r = 2'b10;
			14'b10000111111011: M1r = 2'b10;
			14'b11000111111011: M1r = 2'b10;
			14'b00010111111011: M1r = 2'b01;
			14'b01010111111011: M1r = 2'b01;
			14'b10010111111011: M1r = 2'b10;
			14'b11010111111011: M1r = 2'b10;
			14'b00100111111011: M1r = 2'b01;
			14'b01100111111011: M1r = 2'b01;
			14'b10100111111011: M1r = 2'b01;
			14'b11100111111011: M1r = 2'b01;
			14'b00110111111011: M1r = 2'b00;
			14'b01110111111011: M1r = 2'b00;
			14'b10110111111011: M1r = 2'b01;
			14'b11110111111011: M1r = 2'b01;
			14'b00001011111011: M1r = 2'b10;
			14'b01001011111011: M1r = 2'b11;
			14'b10001011111011: M1r = 2'b11;
			14'b11001011111011: M1r = 2'b11;
			14'b00011011111011: M1r = 2'b10;
			14'b01011011111011: M1r = 2'b10;
			14'b10011011111011: M1r = 2'b10;
			14'b11011011111011: M1r = 2'b10;
			14'b00101011111011: M1r = 2'b10;
			14'b01101011111011: M1r = 2'b10;
			14'b10101011111011: M1r = 2'b10;
			14'b11101011111011: M1r = 2'b10;
			14'b00111011111011: M1r = 2'b01;
			14'b01111011111011: M1r = 2'b01;
			14'b10111011111011: M1r = 2'b01;
			14'b11111011111011: M1r = 2'b10;
			14'b00001111111011: M1r = 2'b11;
			14'b01001111111011: M1r = 2'b11;
			14'b10001111111011: M1r = 2'b11;
			14'b11001111111011: M1r = 2'b11;
			14'b00011111111011: M1r = 2'b11;
			14'b01011111111011: M1r = 2'b11;
			14'b10011111111011: M1r = 2'b11;
			14'b11011111111011: M1r = 2'b11;
			14'b00101111111011: M1r = 2'b10;
			14'b01101111111011: M1r = 2'b10;
			14'b10101111111011: M1r = 2'b11;
			14'b11101111111011: M1r = 2'b11;
			14'b00111111111011: M1r = 2'b10;
			14'b01111111111011: M1r = 2'b10;
			14'b10111111111011: M1r = 2'b10;
			14'b11111111111011: M1r = 2'b10;
			14'b00000000001111: M1r = 2'b00;
			14'b01000000001111: M1r = 2'b00;
			14'b10000000001111: M1r = 2'b00;
			14'b11000000001111: M1r = 2'b00;
			14'b00010000001111: M1r = 2'b00;
			14'b01010000001111: M1r = 2'b00;
			14'b10010000001111: M1r = 2'b00;
			14'b11010000001111: M1r = 2'b00;
			14'b00100000001111: M1r = 2'b00;
			14'b01100000001111: M1r = 2'b00;
			14'b10100000001111: M1r = 2'b00;
			14'b11100000001111: M1r = 2'b00;
			14'b00110000001111: M1r = 2'b00;
			14'b01110000001111: M1r = 2'b00;
			14'b10110000001111: M1r = 2'b00;
			14'b11110000001111: M1r = 2'b00;
			14'b00000100001111: M1r = 2'b00;
			14'b01000100001111: M1r = 2'b01;
			14'b10000100001111: M1r = 2'b01;
			14'b11000100001111: M1r = 2'b01;
			14'b00010100001111: M1r = 2'b00;
			14'b01010100001111: M1r = 2'b00;
			14'b10010100001111: M1r = 2'b00;
			14'b11010100001111: M1r = 2'b00;
			14'b00100100001111: M1r = 2'b00;
			14'b01100100001111: M1r = 2'b00;
			14'b10100100001111: M1r = 2'b00;
			14'b11100100001111: M1r = 2'b00;
			14'b00110100001111: M1r = 2'b00;
			14'b01110100001111: M1r = 2'b00;
			14'b10110100001111: M1r = 2'b00;
			14'b11110100001111: M1r = 2'b00;
			14'b00001000001111: M1r = 2'b01;
			14'b01001000001111: M1r = 2'b01;
			14'b10001000001111: M1r = 2'b10;
			14'b11001000001111: M1r = 2'b10;
			14'b00011000001111: M1r = 2'b01;
			14'b01011000001111: M1r = 2'b01;
			14'b10011000001111: M1r = 2'b01;
			14'b11011000001111: M1r = 2'b01;
			14'b00101000001111: M1r = 2'b00;
			14'b01101000001111: M1r = 2'b00;
			14'b10101000001111: M1r = 2'b01;
			14'b11101000001111: M1r = 2'b01;
			14'b00111000001111: M1r = 2'b00;
			14'b01111000001111: M1r = 2'b00;
			14'b10111000001111: M1r = 2'b00;
			14'b11111000001111: M1r = 2'b00;
			14'b00001100001111: M1r = 2'b10;
			14'b01001100001111: M1r = 2'b10;
			14'b10001100001111: M1r = 2'b10;
			14'b11001100001111: M1r = 2'b10;
			14'b00011100001111: M1r = 2'b01;
			14'b01011100001111: M1r = 2'b10;
			14'b10011100001111: M1r = 2'b10;
			14'b11011100001111: M1r = 2'b10;
			14'b00101100001111: M1r = 2'b01;
			14'b01101100001111: M1r = 2'b01;
			14'b10101100001111: M1r = 2'b01;
			14'b11101100001111: M1r = 2'b01;
			14'b00111100001111: M1r = 2'b01;
			14'b01111100001111: M1r = 2'b01;
			14'b10111100001111: M1r = 2'b01;
			14'b11111100001111: M1r = 2'b01;
			14'b00000001001111: M1r = 2'b00;
			14'b01000001001111: M1r = 2'b00;
			14'b10000001001111: M1r = 2'b00;
			14'b11000001001111: M1r = 2'b00;
			14'b00010001001111: M1r = 2'b00;
			14'b01010001001111: M1r = 2'b00;
			14'b10010001001111: M1r = 2'b00;
			14'b11010001001111: M1r = 2'b00;
			14'b00100001001111: M1r = 2'b00;
			14'b01100001001111: M1r = 2'b00;
			14'b10100001001111: M1r = 2'b00;
			14'b11100001001111: M1r = 2'b00;
			14'b00110001001111: M1r = 2'b00;
			14'b01110001001111: M1r = 2'b00;
			14'b10110001001111: M1r = 2'b00;
			14'b11110001001111: M1r = 2'b00;
			14'b00000101001111: M1r = 2'b00;
			14'b01000101001111: M1r = 2'b00;
			14'b10000101001111: M1r = 2'b00;
			14'b11000101001111: M1r = 2'b01;
			14'b00010101001111: M1r = 2'b00;
			14'b01010101001111: M1r = 2'b00;
			14'b10010101001111: M1r = 2'b00;
			14'b11010101001111: M1r = 2'b00;
			14'b00100101001111: M1r = 2'b00;
			14'b01100101001111: M1r = 2'b00;
			14'b10100101001111: M1r = 2'b00;
			14'b11100101001111: M1r = 2'b00;
			14'b00110101001111: M1r = 2'b00;
			14'b01110101001111: M1r = 2'b00;
			14'b10110101001111: M1r = 2'b00;
			14'b11110101001111: M1r = 2'b00;
			14'b00001001001111: M1r = 2'b01;
			14'b01001001001111: M1r = 2'b01;
			14'b10001001001111: M1r = 2'b01;
			14'b11001001001111: M1r = 2'b01;
			14'b00011001001111: M1r = 2'b00;
			14'b01011001001111: M1r = 2'b01;
			14'b10011001001111: M1r = 2'b01;
			14'b11011001001111: M1r = 2'b01;
			14'b00101001001111: M1r = 2'b00;
			14'b01101001001111: M1r = 2'b00;
			14'b10101001001111: M1r = 2'b00;
			14'b11101001001111: M1r = 2'b00;
			14'b00111001001111: M1r = 2'b00;
			14'b01111001001111: M1r = 2'b00;
			14'b10111001001111: M1r = 2'b00;
			14'b11111001001111: M1r = 2'b00;
			14'b00001101001111: M1r = 2'b10;
			14'b01001101001111: M1r = 2'b10;
			14'b10001101001111: M1r = 2'b10;
			14'b11001101001111: M1r = 2'b10;
			14'b00011101001111: M1r = 2'b01;
			14'b01011101001111: M1r = 2'b01;
			14'b10011101001111: M1r = 2'b10;
			14'b11011101001111: M1r = 2'b10;
			14'b00101101001111: M1r = 2'b01;
			14'b01101101001111: M1r = 2'b01;
			14'b10101101001111: M1r = 2'b01;
			14'b11101101001111: M1r = 2'b01;
			14'b00111101001111: M1r = 2'b00;
			14'b01111101001111: M1r = 2'b00;
			14'b10111101001111: M1r = 2'b01;
			14'b11111101001111: M1r = 2'b01;
			14'b00000010001111: M1r = 2'b00;
			14'b01000010001111: M1r = 2'b00;
			14'b10000010001111: M1r = 2'b00;
			14'b11000010001111: M1r = 2'b00;
			14'b00010010001111: M1r = 2'b00;
			14'b01010010001111: M1r = 2'b00;
			14'b10010010001111: M1r = 2'b00;
			14'b11010010001111: M1r = 2'b00;
			14'b00100010001111: M1r = 2'b00;
			14'b01100010001111: M1r = 2'b00;
			14'b10100010001111: M1r = 2'b00;
			14'b11100010001111: M1r = 2'b00;
			14'b00110010001111: M1r = 2'b00;
			14'b01110010001111: M1r = 2'b00;
			14'b10110010001111: M1r = 2'b00;
			14'b11110010001111: M1r = 2'b00;
			14'b00000110001111: M1r = 2'b00;
			14'b01000110001111: M1r = 2'b00;
			14'b10000110001111: M1r = 2'b00;
			14'b11000110001111: M1r = 2'b00;
			14'b00010110001111: M1r = 2'b00;
			14'b01010110001111: M1r = 2'b00;
			14'b10010110001111: M1r = 2'b00;
			14'b11010110001111: M1r = 2'b00;
			14'b00100110001111: M1r = 2'b00;
			14'b01100110001111: M1r = 2'b00;
			14'b10100110001111: M1r = 2'b00;
			14'b11100110001111: M1r = 2'b00;
			14'b00110110001111: M1r = 2'b00;
			14'b01110110001111: M1r = 2'b00;
			14'b10110110001111: M1r = 2'b00;
			14'b11110110001111: M1r = 2'b00;
			14'b00001010001111: M1r = 2'b01;
			14'b01001010001111: M1r = 2'b01;
			14'b10001010001111: M1r = 2'b01;
			14'b11001010001111: M1r = 2'b01;
			14'b00011010001111: M1r = 2'b00;
			14'b01011010001111: M1r = 2'b00;
			14'b10011010001111: M1r = 2'b00;
			14'b11011010001111: M1r = 2'b01;
			14'b00101010001111: M1r = 2'b00;
			14'b01101010001111: M1r = 2'b00;
			14'b10101010001111: M1r = 2'b00;
			14'b11101010001111: M1r = 2'b00;
			14'b00111010001111: M1r = 2'b00;
			14'b01111010001111: M1r = 2'b00;
			14'b10111010001111: M1r = 2'b00;
			14'b11111010001111: M1r = 2'b00;
			14'b00001110001111: M1r = 2'b01;
			14'b01001110001111: M1r = 2'b10;
			14'b10001110001111: M1r = 2'b10;
			14'b11001110001111: M1r = 2'b10;
			14'b00011110001111: M1r = 2'b01;
			14'b01011110001111: M1r = 2'b01;
			14'b10011110001111: M1r = 2'b01;
			14'b11011110001111: M1r = 2'b01;
			14'b00101110001111: M1r = 2'b00;
			14'b01101110001111: M1r = 2'b01;
			14'b10101110001111: M1r = 2'b01;
			14'b11101110001111: M1r = 2'b01;
			14'b00111110001111: M1r = 2'b00;
			14'b01111110001111: M1r = 2'b00;
			14'b10111110001111: M1r = 2'b00;
			14'b11111110001111: M1r = 2'b00;
			14'b00000011001111: M1r = 2'b00;
			14'b01000011001111: M1r = 2'b00;
			14'b10000011001111: M1r = 2'b00;
			14'b11000011001111: M1r = 2'b00;
			14'b00010011001111: M1r = 2'b00;
			14'b01010011001111: M1r = 2'b00;
			14'b10010011001111: M1r = 2'b00;
			14'b11010011001111: M1r = 2'b00;
			14'b00100011001111: M1r = 2'b00;
			14'b01100011001111: M1r = 2'b00;
			14'b10100011001111: M1r = 2'b00;
			14'b11100011001111: M1r = 2'b00;
			14'b00110011001111: M1r = 2'b00;
			14'b01110011001111: M1r = 2'b00;
			14'b10110011001111: M1r = 2'b00;
			14'b11110011001111: M1r = 2'b00;
			14'b00000111001111: M1r = 2'b00;
			14'b01000111001111: M1r = 2'b00;
			14'b10000111001111: M1r = 2'b00;
			14'b11000111001111: M1r = 2'b00;
			14'b00010111001111: M1r = 2'b00;
			14'b01010111001111: M1r = 2'b00;
			14'b10010111001111: M1r = 2'b00;
			14'b11010111001111: M1r = 2'b00;
			14'b00100111001111: M1r = 2'b00;
			14'b01100111001111: M1r = 2'b00;
			14'b10100111001111: M1r = 2'b00;
			14'b11100111001111: M1r = 2'b00;
			14'b00110111001111: M1r = 2'b00;
			14'b01110111001111: M1r = 2'b00;
			14'b10110111001111: M1r = 2'b00;
			14'b11110111001111: M1r = 2'b00;
			14'b00001011001111: M1r = 2'b00;
			14'b01001011001111: M1r = 2'b01;
			14'b10001011001111: M1r = 2'b01;
			14'b11001011001111: M1r = 2'b01;
			14'b00011011001111: M1r = 2'b00;
			14'b01011011001111: M1r = 2'b00;
			14'b10011011001111: M1r = 2'b00;
			14'b11011011001111: M1r = 2'b00;
			14'b00101011001111: M1r = 2'b00;
			14'b01101011001111: M1r = 2'b00;
			14'b10101011001111: M1r = 2'b00;
			14'b11101011001111: M1r = 2'b00;
			14'b00111011001111: M1r = 2'b00;
			14'b01111011001111: M1r = 2'b00;
			14'b10111011001111: M1r = 2'b00;
			14'b11111011001111: M1r = 2'b00;
			14'b00001111001111: M1r = 2'b01;
			14'b01001111001111: M1r = 2'b01;
			14'b10001111001111: M1r = 2'b01;
			14'b11001111001111: M1r = 2'b10;
			14'b00011111001111: M1r = 2'b01;
			14'b01011111001111: M1r = 2'b01;
			14'b10011111001111: M1r = 2'b01;
			14'b11011111001111: M1r = 2'b01;
			14'b00101111001111: M1r = 2'b00;
			14'b01101111001111: M1r = 2'b00;
			14'b10101111001111: M1r = 2'b00;
			14'b11101111001111: M1r = 2'b01;
			14'b00111111001111: M1r = 2'b00;
			14'b01111111001111: M1r = 2'b00;
			14'b10111111001111: M1r = 2'b00;
			14'b11111111001111: M1r = 2'b00;
			14'b00000000011111: M1r = 2'b00;
			14'b01000000011111: M1r = 2'b00;
			14'b10000000011111: M1r = 2'b00;
			14'b11000000011111: M1r = 2'b01;
			14'b00010000011111: M1r = 2'b00;
			14'b01010000011111: M1r = 2'b00;
			14'b10010000011111: M1r = 2'b00;
			14'b11010000011111: M1r = 2'b00;
			14'b00100000011111: M1r = 2'b00;
			14'b01100000011111: M1r = 2'b00;
			14'b10100000011111: M1r = 2'b00;
			14'b11100000011111: M1r = 2'b00;
			14'b00110000011111: M1r = 2'b00;
			14'b01110000011111: M1r = 2'b00;
			14'b10110000011111: M1r = 2'b00;
			14'b11110000011111: M1r = 2'b00;
			14'b00000100011111: M1r = 2'b01;
			14'b01000100011111: M1r = 2'b01;
			14'b10000100011111: M1r = 2'b01;
			14'b11000100011111: M1r = 2'b01;
			14'b00010100011111: M1r = 2'b00;
			14'b01010100011111: M1r = 2'b01;
			14'b10010100011111: M1r = 2'b01;
			14'b11010100011111: M1r = 2'b01;
			14'b00100100011111: M1r = 2'b00;
			14'b01100100011111: M1r = 2'b00;
			14'b10100100011111: M1r = 2'b00;
			14'b11100100011111: M1r = 2'b00;
			14'b00110100011111: M1r = 2'b00;
			14'b01110100011111: M1r = 2'b00;
			14'b10110100011111: M1r = 2'b00;
			14'b11110100011111: M1r = 2'b00;
			14'b00001000011111: M1r = 2'b10;
			14'b01001000011111: M1r = 2'b10;
			14'b10001000011111: M1r = 2'b10;
			14'b11001000011111: M1r = 2'b10;
			14'b00011000011111: M1r = 2'b01;
			14'b01011000011111: M1r = 2'b01;
			14'b10011000011111: M1r = 2'b01;
			14'b11011000011111: M1r = 2'b10;
			14'b00101000011111: M1r = 2'b01;
			14'b01101000011111: M1r = 2'b01;
			14'b10101000011111: M1r = 2'b01;
			14'b11101000011111: M1r = 2'b01;
			14'b00111000011111: M1r = 2'b00;
			14'b01111000011111: M1r = 2'b00;
			14'b10111000011111: M1r = 2'b01;
			14'b11111000011111: M1r = 2'b01;
			14'b00001100011111: M1r = 2'b10;
			14'b01001100011111: M1r = 2'b11;
			14'b10001100011111: M1r = 2'b11;
			14'b11001100011111: M1r = 2'b11;
			14'b00011100011111: M1r = 2'b10;
			14'b01011100011111: M1r = 2'b10;
			14'b10011100011111: M1r = 2'b10;
			14'b11011100011111: M1r = 2'b10;
			14'b00101100011111: M1r = 2'b01;
			14'b01101100011111: M1r = 2'b10;
			14'b10101100011111: M1r = 2'b10;
			14'b11101100011111: M1r = 2'b10;
			14'b00111100011111: M1r = 2'b01;
			14'b01111100011111: M1r = 2'b01;
			14'b10111100011111: M1r = 2'b01;
			14'b11111100011111: M1r = 2'b01;
			14'b00000001011111: M1r = 2'b00;
			14'b01000001011111: M1r = 2'b00;
			14'b10000001011111: M1r = 2'b00;
			14'b11000001011111: M1r = 2'b00;
			14'b00010001011111: M1r = 2'b00;
			14'b01010001011111: M1r = 2'b00;
			14'b10010001011111: M1r = 2'b00;
			14'b11010001011111: M1r = 2'b00;
			14'b00100001011111: M1r = 2'b00;
			14'b01100001011111: M1r = 2'b00;
			14'b10100001011111: M1r = 2'b00;
			14'b11100001011111: M1r = 2'b00;
			14'b00110001011111: M1r = 2'b00;
			14'b01110001011111: M1r = 2'b00;
			14'b10110001011111: M1r = 2'b00;
			14'b11110001011111: M1r = 2'b00;
			14'b00000101011111: M1r = 2'b01;
			14'b01000101011111: M1r = 2'b01;
			14'b10000101011111: M1r = 2'b01;
			14'b11000101011111: M1r = 2'b01;
			14'b00010101011111: M1r = 2'b00;
			14'b01010101011111: M1r = 2'b00;
			14'b10010101011111: M1r = 2'b00;
			14'b11010101011111: M1r = 2'b01;
			14'b00100101011111: M1r = 2'b00;
			14'b01100101011111: M1r = 2'b00;
			14'b10100101011111: M1r = 2'b00;
			14'b11100101011111: M1r = 2'b00;
			14'b00110101011111: M1r = 2'b00;
			14'b01110101011111: M1r = 2'b00;
			14'b10110101011111: M1r = 2'b00;
			14'b11110101011111: M1r = 2'b00;
			14'b00001001011111: M1r = 2'b01;
			14'b01001001011111: M1r = 2'b10;
			14'b10001001011111: M1r = 2'b10;
			14'b11001001011111: M1r = 2'b10;
			14'b00011001011111: M1r = 2'b01;
			14'b01011001011111: M1r = 2'b01;
			14'b10011001011111: M1r = 2'b01;
			14'b11011001011111: M1r = 2'b01;
			14'b00101001011111: M1r = 2'b00;
			14'b01101001011111: M1r = 2'b01;
			14'b10101001011111: M1r = 2'b01;
			14'b11101001011111: M1r = 2'b01;
			14'b00111001011111: M1r = 2'b00;
			14'b01111001011111: M1r = 2'b00;
			14'b10111001011111: M1r = 2'b00;
			14'b11111001011111: M1r = 2'b00;
			14'b00001101011111: M1r = 2'b10;
			14'b01001101011111: M1r = 2'b10;
			14'b10001101011111: M1r = 2'b10;
			14'b11001101011111: M1r = 2'b11;
			14'b00011101011111: M1r = 2'b10;
			14'b01011101011111: M1r = 2'b10;
			14'b10011101011111: M1r = 2'b10;
			14'b11011101011111: M1r = 2'b10;
			14'b00101101011111: M1r = 2'b01;
			14'b01101101011111: M1r = 2'b01;
			14'b10101101011111: M1r = 2'b01;
			14'b11101101011111: M1r = 2'b10;
			14'b00111101011111: M1r = 2'b01;
			14'b01111101011111: M1r = 2'b01;
			14'b10111101011111: M1r = 2'b01;
			14'b11111101011111: M1r = 2'b01;
			14'b00000010011111: M1r = 2'b00;
			14'b01000010011111: M1r = 2'b00;
			14'b10000010011111: M1r = 2'b00;
			14'b11000010011111: M1r = 2'b00;
			14'b00010010011111: M1r = 2'b00;
			14'b01010010011111: M1r = 2'b00;
			14'b10010010011111: M1r = 2'b00;
			14'b11010010011111: M1r = 2'b00;
			14'b00100010011111: M1r = 2'b00;
			14'b01100010011111: M1r = 2'b00;
			14'b10100010011111: M1r = 2'b00;
			14'b11100010011111: M1r = 2'b00;
			14'b00110010011111: M1r = 2'b00;
			14'b01110010011111: M1r = 2'b00;
			14'b10110010011111: M1r = 2'b00;
			14'b11110010011111: M1r = 2'b00;
			14'b00000110011111: M1r = 2'b00;
			14'b01000110011111: M1r = 2'b00;
			14'b10000110011111: M1r = 2'b01;
			14'b11000110011111: M1r = 2'b01;
			14'b00010110011111: M1r = 2'b00;
			14'b01010110011111: M1r = 2'b00;
			14'b10010110011111: M1r = 2'b00;
			14'b11010110011111: M1r = 2'b00;
			14'b00100110011111: M1r = 2'b00;
			14'b01100110011111: M1r = 2'b00;
			14'b10100110011111: M1r = 2'b00;
			14'b11100110011111: M1r = 2'b00;
			14'b00110110011111: M1r = 2'b00;
			14'b01110110011111: M1r = 2'b00;
			14'b10110110011111: M1r = 2'b00;
			14'b11110110011111: M1r = 2'b00;
			14'b00001010011111: M1r = 2'b01;
			14'b01001010011111: M1r = 2'b01;
			14'b10001010011111: M1r = 2'b01;
			14'b11001010011111: M1r = 2'b10;
			14'b00011010011111: M1r = 2'b01;
			14'b01011010011111: M1r = 2'b01;
			14'b10011010011111: M1r = 2'b01;
			14'b11011010011111: M1r = 2'b01;
			14'b00101010011111: M1r = 2'b00;
			14'b01101010011111: M1r = 2'b00;
			14'b10101010011111: M1r = 2'b00;
			14'b11101010011111: M1r = 2'b01;
			14'b00111010011111: M1r = 2'b00;
			14'b01111010011111: M1r = 2'b00;
			14'b10111010011111: M1r = 2'b00;
			14'b11111010011111: M1r = 2'b00;
			14'b00001110011111: M1r = 2'b10;
			14'b01001110011111: M1r = 2'b10;
			14'b10001110011111: M1r = 2'b10;
			14'b11001110011111: M1r = 2'b10;
			14'b00011110011111: M1r = 2'b01;
			14'b01011110011111: M1r = 2'b10;
			14'b10011110011111: M1r = 2'b10;
			14'b11011110011111: M1r = 2'b10;
			14'b00101110011111: M1r = 2'b01;
			14'b01101110011111: M1r = 2'b01;
			14'b10101110011111: M1r = 2'b01;
			14'b11101110011111: M1r = 2'b01;
			14'b00111110011111: M1r = 2'b00;
			14'b01111110011111: M1r = 2'b01;
			14'b10111110011111: M1r = 2'b01;
			14'b11111110011111: M1r = 2'b01;
			14'b00000011011111: M1r = 2'b00;
			14'b01000011011111: M1r = 2'b00;
			14'b10000011011111: M1r = 2'b00;
			14'b11000011011111: M1r = 2'b00;
			14'b00010011011111: M1r = 2'b00;
			14'b01010011011111: M1r = 2'b00;
			14'b10010011011111: M1r = 2'b00;
			14'b11010011011111: M1r = 2'b00;
			14'b00100011011111: M1r = 2'b00;
			14'b01100011011111: M1r = 2'b00;
			14'b10100011011111: M1r = 2'b00;
			14'b11100011011111: M1r = 2'b00;
			14'b00110011011111: M1r = 2'b00;
			14'b01110011011111: M1r = 2'b00;
			14'b10110011011111: M1r = 2'b00;
			14'b11110011011111: M1r = 2'b00;
			14'b00000111011111: M1r = 2'b00;
			14'b01000111011111: M1r = 2'b00;
			14'b10000111011111: M1r = 2'b00;
			14'b11000111011111: M1r = 2'b01;
			14'b00010111011111: M1r = 2'b00;
			14'b01010111011111: M1r = 2'b00;
			14'b10010111011111: M1r = 2'b00;
			14'b11010111011111: M1r = 2'b00;
			14'b00100111011111: M1r = 2'b00;
			14'b01100111011111: M1r = 2'b00;
			14'b10100111011111: M1r = 2'b00;
			14'b11100111011111: M1r = 2'b00;
			14'b00110111011111: M1r = 2'b00;
			14'b01110111011111: M1r = 2'b00;
			14'b10110111011111: M1r = 2'b00;
			14'b11110111011111: M1r = 2'b00;
			14'b00001011011111: M1r = 2'b01;
			14'b01001011011111: M1r = 2'b01;
			14'b10001011011111: M1r = 2'b01;
			14'b11001011011111: M1r = 2'b01;
			14'b00011011011111: M1r = 2'b00;
			14'b01011011011111: M1r = 2'b00;
			14'b10011011011111: M1r = 2'b01;
			14'b11011011011111: M1r = 2'b01;
			14'b00101011011111: M1r = 2'b00;
			14'b01101011011111: M1r = 2'b00;
			14'b10101011011111: M1r = 2'b00;
			14'b11101011011111: M1r = 2'b00;
			14'b00111011011111: M1r = 2'b00;
			14'b01111011011111: M1r = 2'b00;
			14'b10111011011111: M1r = 2'b00;
			14'b11111011011111: M1r = 2'b00;
			14'b00001111011111: M1r = 2'b10;
			14'b01001111011111: M1r = 2'b10;
			14'b10001111011111: M1r = 2'b10;
			14'b11001111011111: M1r = 2'b10;
			14'b00011111011111: M1r = 2'b01;
			14'b01011111011111: M1r = 2'b01;
			14'b10011111011111: M1r = 2'b01;
			14'b11011111011111: M1r = 2'b10;
			14'b00101111011111: M1r = 2'b01;
			14'b01101111011111: M1r = 2'b01;
			14'b10101111011111: M1r = 2'b01;
			14'b11101111011111: M1r = 2'b01;
			14'b00111111011111: M1r = 2'b00;
			14'b01111111011111: M1r = 2'b00;
			14'b10111111011111: M1r = 2'b00;
			14'b11111111011111: M1r = 2'b01;
			14'b00000000101111: M1r = 2'b01;
			14'b01000000101111: M1r = 2'b01;
			14'b10000000101111: M1r = 2'b01;
			14'b11000000101111: M1r = 2'b01;
			14'b00010000101111: M1r = 2'b00;
			14'b01010000101111: M1r = 2'b00;
			14'b10010000101111: M1r = 2'b00;
			14'b11010000101111: M1r = 2'b01;
			14'b00100000101111: M1r = 2'b00;
			14'b01100000101111: M1r = 2'b00;
			14'b10100000101111: M1r = 2'b00;
			14'b11100000101111: M1r = 2'b00;
			14'b00110000101111: M1r = 2'b00;
			14'b01110000101111: M1r = 2'b00;
			14'b10110000101111: M1r = 2'b00;
			14'b11110000101111: M1r = 2'b00;
			14'b00000100101111: M1r = 2'b01;
			14'b01000100101111: M1r = 2'b01;
			14'b10000100101111: M1r = 2'b10;
			14'b11000100101111: M1r = 2'b10;
			14'b00010100101111: M1r = 2'b01;
			14'b01010100101111: M1r = 2'b01;
			14'b10010100101111: M1r = 2'b01;
			14'b11010100101111: M1r = 2'b01;
			14'b00100100101111: M1r = 2'b00;
			14'b01100100101111: M1r = 2'b01;
			14'b10100100101111: M1r = 2'b01;
			14'b11100100101111: M1r = 2'b01;
			14'b00110100101111: M1r = 2'b00;
			14'b01110100101111: M1r = 2'b00;
			14'b10110100101111: M1r = 2'b00;
			14'b11110100101111: M1r = 2'b00;
			14'b00001000101111: M1r = 2'b10;
			14'b01001000101111: M1r = 2'b10;
			14'b10001000101111: M1r = 2'b10;
			14'b11001000101111: M1r = 2'b11;
			14'b00011000101111: M1r = 2'b10;
			14'b01011000101111: M1r = 2'b10;
			14'b10011000101111: M1r = 2'b10;
			14'b11011000101111: M1r = 2'b10;
			14'b00101000101111: M1r = 2'b01;
			14'b01101000101111: M1r = 2'b01;
			14'b10101000101111: M1r = 2'b01;
			14'b11101000101111: M1r = 2'b10;
			14'b00111000101111: M1r = 2'b01;
			14'b01111000101111: M1r = 2'b01;
			14'b10111000101111: M1r = 2'b01;
			14'b11111000101111: M1r = 2'b01;
			14'b00001100101111: M1r = 2'b11;
			14'b01001100101111: M1r = 2'b11;
			14'b10001100101111: M1r = 2'b11;
			14'b11001100101111: M1r = 2'b11;
			14'b00011100101111: M1r = 2'b10;
			14'b01011100101111: M1r = 2'b11;
			14'b10011100101111: M1r = 2'b11;
			14'b11011100101111: M1r = 2'b11;
			14'b00101100101111: M1r = 2'b10;
			14'b01101100101111: M1r = 2'b10;
			14'b10101100101111: M1r = 2'b10;
			14'b11101100101111: M1r = 2'b10;
			14'b00111100101111: M1r = 2'b01;
			14'b01111100101111: M1r = 2'b10;
			14'b10111100101111: M1r = 2'b10;
			14'b11111100101111: M1r = 2'b10;
			14'b00000001101111: M1r = 2'b00;
			14'b01000001101111: M1r = 2'b00;
			14'b10000001101111: M1r = 2'b01;
			14'b11000001101111: M1r = 2'b01;
			14'b00010001101111: M1r = 2'b00;
			14'b01010001101111: M1r = 2'b00;
			14'b10010001101111: M1r = 2'b00;
			14'b11010001101111: M1r = 2'b00;
			14'b00100001101111: M1r = 2'b00;
			14'b01100001101111: M1r = 2'b00;
			14'b10100001101111: M1r = 2'b00;
			14'b11100001101111: M1r = 2'b00;
			14'b00110001101111: M1r = 2'b00;
			14'b01110001101111: M1r = 2'b00;
			14'b10110001101111: M1r = 2'b00;
			14'b11110001101111: M1r = 2'b00;
			14'b00000101101111: M1r = 2'b01;
			14'b01000101101111: M1r = 2'b01;
			14'b10000101101111: M1r = 2'b01;
			14'b11000101101111: M1r = 2'b10;
			14'b00010101101111: M1r = 2'b01;
			14'b01010101101111: M1r = 2'b01;
			14'b10010101101111: M1r = 2'b01;
			14'b11010101101111: M1r = 2'b01;
			14'b00100101101111: M1r = 2'b00;
			14'b01100101101111: M1r = 2'b00;
			14'b10100101101111: M1r = 2'b00;
			14'b11100101101111: M1r = 2'b01;
			14'b00110101101111: M1r = 2'b00;
			14'b01110101101111: M1r = 2'b00;
			14'b10110101101111: M1r = 2'b00;
			14'b11110101101111: M1r = 2'b00;
			14'b00001001101111: M1r = 2'b10;
			14'b01001001101111: M1r = 2'b10;
			14'b10001001101111: M1r = 2'b10;
			14'b11001001101111: M1r = 2'b10;
			14'b00011001101111: M1r = 2'b01;
			14'b01011001101111: M1r = 2'b01;
			14'b10011001101111: M1r = 2'b10;
			14'b11011001101111: M1r = 2'b10;
			14'b00101001101111: M1r = 2'b01;
			14'b01101001101111: M1r = 2'b01;
			14'b10101001101111: M1r = 2'b01;
			14'b11101001101111: M1r = 2'b01;
			14'b00111001101111: M1r = 2'b00;
			14'b01111001101111: M1r = 2'b01;
			14'b10111001101111: M1r = 2'b01;
			14'b11111001101111: M1r = 2'b01;
			14'b00001101101111: M1r = 2'b11;
			14'b01001101101111: M1r = 2'b11;
			14'b10001101101111: M1r = 2'b11;
			14'b11001101101111: M1r = 2'b11;
			14'b00011101101111: M1r = 2'b10;
			14'b01011101101111: M1r = 2'b10;
			14'b10011101101111: M1r = 2'b10;
			14'b11011101101111: M1r = 2'b11;
			14'b00101101101111: M1r = 2'b10;
			14'b01101101101111: M1r = 2'b10;
			14'b10101101101111: M1r = 2'b10;
			14'b11101101101111: M1r = 2'b10;
			14'b00111101101111: M1r = 2'b01;
			14'b01111101101111: M1r = 2'b01;
			14'b10111101101111: M1r = 2'b01;
			14'b11111101101111: M1r = 2'b10;
			14'b00000010101111: M1r = 2'b00;
			14'b01000010101111: M1r = 2'b00;
			14'b10000010101111: M1r = 2'b00;
			14'b11000010101111: M1r = 2'b00;
			14'b00010010101111: M1r = 2'b00;
			14'b01010010101111: M1r = 2'b00;
			14'b10010010101111: M1r = 2'b00;
			14'b11010010101111: M1r = 2'b00;
			14'b00100010101111: M1r = 2'b00;
			14'b01100010101111: M1r = 2'b00;
			14'b10100010101111: M1r = 2'b00;
			14'b11100010101111: M1r = 2'b00;
			14'b00110010101111: M1r = 2'b00;
			14'b01110010101111: M1r = 2'b00;
			14'b10110010101111: M1r = 2'b00;
			14'b11110010101111: M1r = 2'b00;
			14'b00000110101111: M1r = 2'b01;
			14'b01000110101111: M1r = 2'b01;
			14'b10000110101111: M1r = 2'b01;
			14'b11000110101111: M1r = 2'b01;
			14'b00010110101111: M1r = 2'b00;
			14'b01010110101111: M1r = 2'b00;
			14'b10010110101111: M1r = 2'b01;
			14'b11010110101111: M1r = 2'b01;
			14'b00100110101111: M1r = 2'b00;
			14'b01100110101111: M1r = 2'b00;
			14'b10100110101111: M1r = 2'b00;
			14'b11100110101111: M1r = 2'b00;
			14'b00110110101111: M1r = 2'b00;
			14'b01110110101111: M1r = 2'b00;
			14'b10110110101111: M1r = 2'b00;
			14'b11110110101111: M1r = 2'b00;
			14'b00001010101111: M1r = 2'b10;
			14'b01001010101111: M1r = 2'b10;
			14'b10001010101111: M1r = 2'b10;
			14'b11001010101111: M1r = 2'b10;
			14'b00011010101111: M1r = 2'b01;
			14'b01011010101111: M1r = 2'b01;
			14'b10011010101111: M1r = 2'b01;
			14'b11011010101111: M1r = 2'b10;
			14'b00101010101111: M1r = 2'b01;
			14'b01101010101111: M1r = 2'b01;
			14'b10101010101111: M1r = 2'b01;
			14'b11101010101111: M1r = 2'b01;
			14'b00111010101111: M1r = 2'b00;
			14'b01111010101111: M1r = 2'b00;
			14'b10111010101111: M1r = 2'b00;
			14'b11111010101111: M1r = 2'b01;
			14'b00001110101111: M1r = 2'b10;
			14'b01001110101111: M1r = 2'b10;
			14'b10001110101111: M1r = 2'b11;
			14'b11001110101111: M1r = 2'b11;
			14'b00011110101111: M1r = 2'b10;
			14'b01011110101111: M1r = 2'b10;
			14'b10011110101111: M1r = 2'b10;
			14'b11011110101111: M1r = 2'b10;
			14'b00101110101111: M1r = 2'b01;
			14'b01101110101111: M1r = 2'b01;
			14'b10101110101111: M1r = 2'b10;
			14'b11101110101111: M1r = 2'b10;
			14'b00111110101111: M1r = 2'b01;
			14'b01111110101111: M1r = 2'b01;
			14'b10111110101111: M1r = 2'b01;
			14'b11111110101111: M1r = 2'b01;
			14'b00000011101111: M1r = 2'b00;
			14'b01000011101111: M1r = 2'b00;
			14'b10000011101111: M1r = 2'b00;
			14'b11000011101111: M1r = 2'b00;
			14'b00010011101111: M1r = 2'b00;
			14'b01010011101111: M1r = 2'b00;
			14'b10010011101111: M1r = 2'b00;
			14'b11010011101111: M1r = 2'b00;
			14'b00100011101111: M1r = 2'b00;
			14'b01100011101111: M1r = 2'b00;
			14'b10100011101111: M1r = 2'b00;
			14'b11100011101111: M1r = 2'b00;
			14'b00110011101111: M1r = 2'b00;
			14'b01110011101111: M1r = 2'b00;
			14'b10110011101111: M1r = 2'b00;
			14'b11110011101111: M1r = 2'b00;
			14'b00000111101111: M1r = 2'b01;
			14'b01000111101111: M1r = 2'b01;
			14'b10000111101111: M1r = 2'b01;
			14'b11000111101111: M1r = 2'b01;
			14'b00010111101111: M1r = 2'b00;
			14'b01010111101111: M1r = 2'b00;
			14'b10010111101111: M1r = 2'b00;
			14'b11010111101111: M1r = 2'b00;
			14'b00100111101111: M1r = 2'b00;
			14'b01100111101111: M1r = 2'b00;
			14'b10100111101111: M1r = 2'b00;
			14'b11100111101111: M1r = 2'b00;
			14'b00110111101111: M1r = 2'b00;
			14'b01110111101111: M1r = 2'b00;
			14'b10110111101111: M1r = 2'b00;
			14'b11110111101111: M1r = 2'b00;
			14'b00001011101111: M1r = 2'b01;
			14'b01001011101111: M1r = 2'b01;
			14'b10001011101111: M1r = 2'b10;
			14'b11001011101111: M1r = 2'b10;
			14'b00011011101111: M1r = 2'b01;
			14'b01011011101111: M1r = 2'b01;
			14'b10011011101111: M1r = 2'b01;
			14'b11011011101111: M1r = 2'b01;
			14'b00101011101111: M1r = 2'b00;
			14'b01101011101111: M1r = 2'b00;
			14'b10101011101111: M1r = 2'b01;
			14'b11101011101111: M1r = 2'b01;
			14'b00111011101111: M1r = 2'b00;
			14'b01111011101111: M1r = 2'b00;
			14'b10111011101111: M1r = 2'b00;
			14'b11111011101111: M1r = 2'b00;
			14'b00001111101111: M1r = 2'b10;
			14'b01001111101111: M1r = 2'b10;
			14'b10001111101111: M1r = 2'b10;
			14'b11001111101111: M1r = 2'b10;
			14'b00011111101111: M1r = 2'b10;
			14'b01011111101111: M1r = 2'b10;
			14'b10011111101111: M1r = 2'b10;
			14'b11011111101111: M1r = 2'b10;
			14'b00101111101111: M1r = 2'b01;
			14'b01101111101111: M1r = 2'b01;
			14'b10101111101111: M1r = 2'b01;
			14'b11101111101111: M1r = 2'b10;
			14'b00111111101111: M1r = 2'b01;
			14'b01111111101111: M1r = 2'b01;
			14'b10111111101111: M1r = 2'b01;
			14'b11111111101111: M1r = 2'b01;
			14'b00000000111111: M1r = 2'b01;
			14'b01000000111111: M1r = 2'b01;
			14'b10000000111111: M1r = 2'b01;
			14'b11000000111111: M1r = 2'b01;
			14'b00010000111111: M1r = 2'b01;
			14'b01010000111111: M1r = 2'b01;
			14'b10010000111111: M1r = 2'b01;
			14'b11010000111111: M1r = 2'b01;
			14'b00100000111111: M1r = 2'b00;
			14'b01100000111111: M1r = 2'b00;
			14'b10100000111111: M1r = 2'b00;
			14'b11100000111111: M1r = 2'b01;
			14'b00110000111111: M1r = 2'b00;
			14'b01110000111111: M1r = 2'b00;
			14'b10110000111111: M1r = 2'b00;
			14'b11110000111111: M1r = 2'b00;
			14'b00000100111111: M1r = 2'b10;
			14'b01000100111111: M1r = 2'b10;
			14'b10000100111111: M1r = 2'b10;
			14'b11000100111111: M1r = 2'b10;
			14'b00010100111111: M1r = 2'b01;
			14'b01010100111111: M1r = 2'b01;
			14'b10010100111111: M1r = 2'b10;
			14'b11010100111111: M1r = 2'b10;
			14'b00100100111111: M1r = 2'b01;
			14'b01100100111111: M1r = 2'b01;
			14'b10100100111111: M1r = 2'b01;
			14'b11100100111111: M1r = 2'b01;
			14'b00110100111111: M1r = 2'b00;
			14'b01110100111111: M1r = 2'b00;
			14'b10110100111111: M1r = 2'b01;
			14'b11110100111111: M1r = 2'b01;
			14'b00001000111111: M1r = 2'b11;
			14'b01001000111111: M1r = 2'b11;
			14'b10001000111111: M1r = 2'b11;
			14'b11001000111111: M1r = 2'b11;
			14'b00011000111111: M1r = 2'b10;
			14'b01011000111111: M1r = 2'b10;
			14'b10011000111111: M1r = 2'b10;
			14'b11011000111111: M1r = 2'b10;
			14'b00101000111111: M1r = 2'b10;
			14'b01101000111111: M1r = 2'b10;
			14'b10101000111111: M1r = 2'b10;
			14'b11101000111111: M1r = 2'b10;
			14'b00111000111111: M1r = 2'b01;
			14'b01111000111111: M1r = 2'b01;
			14'b10111000111111: M1r = 2'b01;
			14'b11111000111111: M1r = 2'b10;
			14'b00001100111111: M1r = 2'b11;
			14'b01001100111111: M1r = 2'b11;
			14'b10001100111111: M1r = 2'b11;
			14'b11001100111111: M1r = 2'b11;
			14'b00011100111111: M1r = 2'b11;
			14'b01011100111111: M1r = 2'b11;
			14'b10011100111111: M1r = 2'b11;
			14'b11011100111111: M1r = 2'b11;
			14'b00101100111111: M1r = 2'b10;
			14'b01101100111111: M1r = 2'b10;
			14'b10101100111111: M1r = 2'b11;
			14'b11101100111111: M1r = 2'b11;
			14'b00111100111111: M1r = 2'b10;
			14'b01111100111111: M1r = 2'b10;
			14'b10111100111111: M1r = 2'b10;
			14'b11111100111111: M1r = 2'b10;
			14'b00000001111111: M1r = 2'b01;
			14'b01000001111111: M1r = 2'b01;
			14'b10000001111111: M1r = 2'b01;
			14'b11000001111111: M1r = 2'b01;
			14'b00010001111111: M1r = 2'b00;
			14'b01010001111111: M1r = 2'b00;
			14'b10010001111111: M1r = 2'b01;
			14'b11010001111111: M1r = 2'b01;
			14'b00100001111111: M1r = 2'b00;
			14'b01100001111111: M1r = 2'b00;
			14'b10100001111111: M1r = 2'b00;
			14'b11100001111111: M1r = 2'b00;
			14'b00110001111111: M1r = 2'b00;
			14'b01110001111111: M1r = 2'b00;
			14'b10110001111111: M1r = 2'b00;
			14'b11110001111111: M1r = 2'b00;
			14'b00000101111111: M1r = 2'b01;
			14'b01000101111111: M1r = 2'b10;
			14'b10000101111111: M1r = 2'b10;
			14'b11000101111111: M1r = 2'b10;
			14'b00010101111111: M1r = 2'b01;
			14'b01010101111111: M1r = 2'b01;
			14'b10010101111111: M1r = 2'b01;
			14'b11010101111111: M1r = 2'b01;
			14'b00100101111111: M1r = 2'b01;
			14'b01100101111111: M1r = 2'b01;
			14'b10100101111111: M1r = 2'b01;
			14'b11100101111111: M1r = 2'b01;
			14'b00110101111111: M1r = 2'b00;
			14'b01110101111111: M1r = 2'b00;
			14'b10110101111111: M1r = 2'b00;
			14'b11110101111111: M1r = 2'b01;
			14'b00001001111111: M1r = 2'b10;
			14'b01001001111111: M1r = 2'b10;
			14'b10001001111111: M1r = 2'b11;
			14'b11001001111111: M1r = 2'b11;
			14'b00011001111111: M1r = 2'b10;
			14'b01011001111111: M1r = 2'b10;
			14'b10011001111111: M1r = 2'b10;
			14'b11011001111111: M1r = 2'b10;
			14'b00101001111111: M1r = 2'b01;
			14'b01101001111111: M1r = 2'b01;
			14'b10101001111111: M1r = 2'b10;
			14'b11101001111111: M1r = 2'b10;
			14'b00111001111111: M1r = 2'b01;
			14'b01111001111111: M1r = 2'b01;
			14'b10111001111111: M1r = 2'b01;
			14'b11111001111111: M1r = 2'b01;
			14'b00001101111111: M1r = 2'b11;
			14'b01001101111111: M1r = 2'b11;
			14'b10001101111111: M1r = 2'b11;
			14'b11001101111111: M1r = 2'b11;
			14'b00011101111111: M1r = 2'b11;
			14'b01011101111111: M1r = 2'b11;
			14'b10011101111111: M1r = 2'b11;
			14'b11011101111111: M1r = 2'b11;
			14'b00101101111111: M1r = 2'b10;
			14'b01101101111111: M1r = 2'b10;
			14'b10101101111111: M1r = 2'b10;
			14'b11101101111111: M1r = 2'b10;
			14'b00111101111111: M1r = 2'b10;
			14'b01111101111111: M1r = 2'b10;
			14'b10111101111111: M1r = 2'b10;
			14'b11111101111111: M1r = 2'b10;
			14'b00000010111111: M1r = 2'b00;
			14'b01000010111111: M1r = 2'b01;
			14'b10000010111111: M1r = 2'b01;
			14'b11000010111111: M1r = 2'b01;
			14'b00010010111111: M1r = 2'b00;
			14'b01010010111111: M1r = 2'b00;
			14'b10010010111111: M1r = 2'b00;
			14'b11010010111111: M1r = 2'b00;
			14'b00100010111111: M1r = 2'b00;
			14'b01100010111111: M1r = 2'b00;
			14'b10100010111111: M1r = 2'b00;
			14'b11100010111111: M1r = 2'b00;
			14'b00110010111111: M1r = 2'b00;
			14'b01110010111111: M1r = 2'b00;
			14'b10110010111111: M1r = 2'b00;
			14'b11110010111111: M1r = 2'b00;
			14'b00000110111111: M1r = 2'b01;
			14'b01000110111111: M1r = 2'b01;
			14'b10000110111111: M1r = 2'b10;
			14'b11000110111111: M1r = 2'b10;
			14'b00010110111111: M1r = 2'b01;
			14'b01010110111111: M1r = 2'b01;
			14'b10010110111111: M1r = 2'b01;
			14'b11010110111111: M1r = 2'b01;
			14'b00100110111111: M1r = 2'b00;
			14'b01100110111111: M1r = 2'b00;
			14'b10100110111111: M1r = 2'b01;
			14'b11100110111111: M1r = 2'b01;
			14'b00110110111111: M1r = 2'b00;
			14'b01110110111111: M1r = 2'b00;
			14'b10110110111111: M1r = 2'b00;
			14'b11110110111111: M1r = 2'b00;
			14'b00001010111111: M1r = 2'b10;
			14'b01001010111111: M1r = 2'b10;
			14'b10001010111111: M1r = 2'b10;
			14'b11001010111111: M1r = 2'b10;
			14'b00011010111111: M1r = 2'b01;
			14'b01011010111111: M1r = 2'b10;
			14'b10011010111111: M1r = 2'b10;
			14'b11011010111111: M1r = 2'b10;
			14'b00101010111111: M1r = 2'b01;
			14'b01101010111111: M1r = 2'b01;
			14'b10101010111111: M1r = 2'b01;
			14'b11101010111111: M1r = 2'b01;
			14'b00111010111111: M1r = 2'b01;
			14'b01111010111111: M1r = 2'b01;
			14'b10111010111111: M1r = 2'b01;
			14'b11111010111111: M1r = 2'b01;
			14'b00001110111111: M1r = 2'b11;
			14'b01001110111111: M1r = 2'b11;
			14'b10001110111111: M1r = 2'b11;
			14'b11001110111111: M1r = 2'b11;
			14'b00011110111111: M1r = 2'b10;
			14'b01011110111111: M1r = 2'b10;
			14'b10011110111111: M1r = 2'b11;
			14'b11011110111111: M1r = 2'b11;
			14'b00101110111111: M1r = 2'b10;
			14'b01101110111111: M1r = 2'b10;
			14'b10101110111111: M1r = 2'b10;
			14'b11101110111111: M1r = 2'b10;
			14'b00111110111111: M1r = 2'b01;
			14'b01111110111111: M1r = 2'b01;
			14'b10111110111111: M1r = 2'b10;
			14'b11111110111111: M1r = 2'b10;
			14'b00000011111111: M1r = 2'b00;
			14'b01000011111111: M1r = 2'b00;
			14'b10000011111111: M1r = 2'b00;
			14'b11000011111111: M1r = 2'b01;
			14'b00010011111111: M1r = 2'b00;
			14'b01010011111111: M1r = 2'b00;
			14'b10010011111111: M1r = 2'b00;
			14'b11010011111111: M1r = 2'b00;
			14'b00100011111111: M1r = 2'b00;
			14'b01100011111111: M1r = 2'b00;
			14'b10100011111111: M1r = 2'b00;
			14'b11100011111111: M1r = 2'b00;
			14'b00110011111111: M1r = 2'b00;
			14'b01110011111111: M1r = 2'b00;
			14'b10110011111111: M1r = 2'b00;
			14'b11110011111111: M1r = 2'b00;
			14'b00000111111111: M1r = 2'b01;
			14'b01000111111111: M1r = 2'b01;
			14'b10000111111111: M1r = 2'b01;
			14'b11000111111111: M1r = 2'b01;
			14'b00010111111111: M1r = 2'b00;
			14'b01010111111111: M1r = 2'b01;
			14'b10010111111111: M1r = 2'b01;
			14'b11010111111111: M1r = 2'b01;
			14'b00100111111111: M1r = 2'b00;
			14'b01100111111111: M1r = 2'b00;
			14'b10100111111111: M1r = 2'b00;
			14'b11100111111111: M1r = 2'b00;
			14'b00110111111111: M1r = 2'b00;
			14'b01110111111111: M1r = 2'b00;
			14'b10110111111111: M1r = 2'b00;
			14'b11110111111111: M1r = 2'b00;
			14'b00001011111111: M1r = 2'b10;
			14'b01001011111111: M1r = 2'b10;
			14'b10001011111111: M1r = 2'b10;
			14'b11001011111111: M1r = 2'b10;
			14'b00011011111111: M1r = 2'b01;
			14'b01011011111111: M1r = 2'b01;
			14'b10011011111111: M1r = 2'b10;
			14'b11011011111111: M1r = 2'b10;
			14'b00101011111111: M1r = 2'b01;
			14'b01101011111111: M1r = 2'b01;
			14'b10101011111111: M1r = 2'b01;
			14'b11101011111111: M1r = 2'b01;
			14'b00111011111111: M1r = 2'b00;
			14'b01111011111111: M1r = 2'b00;
			14'b10111011111111: M1r = 2'b01;
			14'b11111011111111: M1r = 2'b01;
			14'b00001111111111: M1r = 2'b10;
			14'b01001111111111: M1r = 2'b11;
			14'b10001111111111: M1r = 2'b11;
			14'b11001111111111: M1r = 2'b11;
			14'b00011111111111: M1r = 2'b10;
			14'b01011111111111: M1r = 2'b10;
			14'b10011111111111: M1r = 2'b10;
			14'b11011111111111: M1r = 2'b10;
			14'b00101111111111: M1r = 2'b01;
			14'b01101111111111: M1r = 2'b10;
			14'b10101111111111: M1r = 2'b10;
			14'b11101111111111: M1r = 2'b10;
			14'b00111111111111: M1r = 2'b01;
			14'b01111111111111: M1r = 2'b01;
			14'b10111111111111: M1r = 2'b01;
			14'b11111111111111: M1r = 2'b01;

		endcase
	end
endmodule
