module layer0_N202 ( input [5:0] M0, output [1:0] M1 );

	(*rom_style = "distributed" *) reg [1:0] M1r;
	assign M1 = M1r;
	always @ (M0) begin
		case (M0)
			6'b000000: M1r = 2'b00;
			6'b100000: M1r = 2'b00;
			6'b010000: M1r = 2'b00;
			6'b110000: M1r = 2'b00;
			6'b001000: M1r = 2'b00;
			6'b101000: M1r = 2'b00;
			6'b011000: M1r = 2'b00;
			6'b111000: M1r = 2'b00;
			6'b000100: M1r = 2'b00;
			6'b100100: M1r = 2'b00;
			6'b010100: M1r = 2'b00;
			6'b110100: M1r = 2'b00;
			6'b001100: M1r = 2'b00;
			6'b101100: M1r = 2'b00;
			6'b011100: M1r = 2'b00;
			6'b111100: M1r = 2'b00;
			6'b000010: M1r = 2'b00;
			6'b100010: M1r = 2'b00;
			6'b010010: M1r = 2'b00;
			6'b110010: M1r = 2'b00;
			6'b001010: M1r = 2'b00;
			6'b101010: M1r = 2'b00;
			6'b011010: M1r = 2'b00;
			6'b111010: M1r = 2'b00;
			6'b000110: M1r = 2'b00;
			6'b100110: M1r = 2'b00;
			6'b010110: M1r = 2'b00;
			6'b110110: M1r = 2'b00;
			6'b001110: M1r = 2'b00;
			6'b101110: M1r = 2'b00;
			6'b011110: M1r = 2'b00;
			6'b111110: M1r = 2'b00;
			6'b000001: M1r = 2'b01;
			6'b100001: M1r = 2'b01;
			6'b010001: M1r = 2'b00;
			6'b110001: M1r = 2'b00;
			6'b001001: M1r = 2'b00;
			6'b101001: M1r = 2'b00;
			6'b011001: M1r = 2'b00;
			6'b111001: M1r = 2'b00;
			6'b000101: M1r = 2'b01;
			6'b100101: M1r = 2'b01;
			6'b010101: M1r = 2'b00;
			6'b110101: M1r = 2'b00;
			6'b001101: M1r = 2'b00;
			6'b101101: M1r = 2'b00;
			6'b011101: M1r = 2'b00;
			6'b111101: M1r = 2'b00;
			6'b000011: M1r = 2'b11;
			6'b100011: M1r = 2'b10;
			6'b010011: M1r = 2'b00;
			6'b110011: M1r = 2'b00;
			6'b001011: M1r = 2'b01;
			6'b101011: M1r = 2'b01;
			6'b011011: M1r = 2'b00;
			6'b111011: M1r = 2'b00;
			6'b000111: M1r = 2'b11;
			6'b100111: M1r = 2'b11;
			6'b010111: M1r = 2'b00;
			6'b110111: M1r = 2'b00;
			6'b001111: M1r = 2'b01;
			6'b101111: M1r = 2'b01;
			6'b011111: M1r = 2'b00;
			6'b111111: M1r = 2'b00;

		endcase
	end
endmodule
