module layer1 (input [511:0] M0, output [171:0] M1);

wire [5:0] layer1_N0_wire = {M0[421], M0[420], M0[65], M0[64], M0[39], M0[38]};
layer1_N0 layer1_N0_inst (.M0(layer1_N0_wire), .M1(M1[1:0]));

wire [5:0] layer1_N1_wire = {M0[451], M0[450], M0[219], M0[218], M0[25], M0[24]};
layer1_N1 layer1_N1_inst (.M0(layer1_N1_wire), .M1(M1[3:2]));

wire [5:0] layer1_N2_wire = {M0[401], M0[400], M0[195], M0[194], M0[181], M0[180]};
layer1_N2 layer1_N2_inst (.M0(layer1_N2_wire), .M1(M1[5:4]));

wire [5:0] layer1_N3_wire = {M0[253], M0[252], M0[159], M0[158], M0[59], M0[58]};
layer1_N3 layer1_N3_inst (.M0(layer1_N3_wire), .M1(M1[7:6]));

wire [5:0] layer1_N4_wire = {M0[335], M0[334], M0[283], M0[282], M0[73], M0[72]};
layer1_N4 layer1_N4_inst (.M0(layer1_N4_wire), .M1(M1[9:8]));

wire [5:0] layer1_N5_wire = {M0[379], M0[378], M0[49], M0[48], M0[41], M0[40]};
layer1_N5 layer1_N5_inst (.M0(layer1_N5_wire), .M1(M1[11:10]));

wire [5:0] layer1_N6_wire = {M0[415], M0[414], M0[229], M0[228], M0[107], M0[106]};
layer1_N6 layer1_N6_inst (.M0(layer1_N6_wire), .M1(M1[13:12]));

wire [5:0] layer1_N7_wire = {M0[203], M0[202], M0[189], M0[188], M0[69], M0[68]};
layer1_N7 layer1_N7_inst (.M0(layer1_N7_wire), .M1(M1[15:14]));

wire [5:0] layer1_N8_wire = {M0[303], M0[302], M0[243], M0[242], M0[173], M0[172]};
layer1_N8 layer1_N8_inst (.M0(layer1_N8_wire), .M1(M1[17:16]));

wire [5:0] layer1_N9_wire = {M0[469], M0[468], M0[431], M0[430], M0[341], M0[340]};
layer1_N9 layer1_N9_inst (.M0(layer1_N9_wire), .M1(M1[19:18]));

wire [5:0] layer1_N10_wire = {M0[415], M0[414], M0[251], M0[250], M0[109], M0[108]};
layer1_N10 layer1_N10_inst (.M0(layer1_N10_wire), .M1(M1[21:20]));

wire [5:0] layer1_N11_wire = {M0[383], M0[382], M0[201], M0[200], M0[159], M0[158]};
layer1_N11 layer1_N11_inst (.M0(layer1_N11_wire), .M1(M1[23:22]));

wire [5:0] layer1_N12_wire = {M0[297], M0[296], M0[287], M0[286], M0[83], M0[82]};
layer1_N12 layer1_N12_inst (.M0(layer1_N12_wire), .M1(M1[25:24]));

wire [5:0] layer1_N13_wire = {M0[505], M0[504], M0[487], M0[486], M0[437], M0[436]};
layer1_N13 layer1_N13_inst (.M0(layer1_N13_wire), .M1(M1[27:26]));

wire [5:0] layer1_N14_wire = {M0[483], M0[482], M0[141], M0[140], M0[87], M0[86]};
layer1_N14 layer1_N14_inst (.M0(layer1_N14_wire), .M1(M1[29:28]));

wire [5:0] layer1_N15_wire = {M0[417], M0[416], M0[225], M0[224], M0[9], M0[8]};
layer1_N15 layer1_N15_inst (.M0(layer1_N15_wire), .M1(M1[31:30]));

wire [5:0] layer1_N16_wire = {M0[187], M0[186], M0[155], M0[154], M0[41], M0[40]};
layer1_N16 layer1_N16_inst (.M0(layer1_N16_wire), .M1(M1[33:32]));

wire [5:0] layer1_N17_wire = {M0[351], M0[350], M0[19], M0[18], M0[15], M0[14]};
layer1_N17 layer1_N17_inst (.M0(layer1_N17_wire), .M1(M1[35:34]));

wire [5:0] layer1_N18_wire = {M0[267], M0[266], M0[221], M0[220], M0[161], M0[160]};
layer1_N18 layer1_N18_inst (.M0(layer1_N18_wire), .M1(M1[37:36]));

wire [5:0] layer1_N19_wire = {M0[189], M0[188], M0[125], M0[124], M0[13], M0[12]};
layer1_N19 layer1_N19_inst (.M0(layer1_N19_wire), .M1(M1[39:38]));

wire [5:0] layer1_N20_wire = {M0[367], M0[366], M0[311], M0[310], M0[69], M0[68]};
layer1_N20 layer1_N20_inst (.M0(layer1_N20_wire), .M1(M1[41:40]));

wire [5:0] layer1_N21_wire = {M0[419], M0[418], M0[139], M0[138], M0[45], M0[44]};
layer1_N21 layer1_N21_inst (.M0(layer1_N21_wire), .M1(M1[43:42]));

wire [5:0] layer1_N22_wire = {M0[473], M0[472], M0[413], M0[412], M0[145], M0[144]};
layer1_N22 layer1_N22_inst (.M0(layer1_N22_wire), .M1(M1[45:44]));

wire [5:0] layer1_N23_wire = {M0[257], M0[256], M0[67], M0[66], M0[15], M0[14]};
layer1_N23 layer1_N23_inst (.M0(layer1_N23_wire), .M1(M1[47:46]));

wire [5:0] layer1_N24_wire = {M0[485], M0[484], M0[303], M0[302], M0[143], M0[142]};
layer1_N24 layer1_N24_inst (.M0(layer1_N24_wire), .M1(M1[49:48]));

wire [5:0] layer1_N25_wire = {M0[497], M0[496], M0[431], M0[430], M0[385], M0[384]};
layer1_N25 layer1_N25_inst (.M0(layer1_N25_wire), .M1(M1[51:50]));

wire [5:0] layer1_N26_wire = {M0[323], M0[322], M0[291], M0[290], M0[233], M0[232]};
layer1_N26 layer1_N26_inst (.M0(layer1_N26_wire), .M1(M1[53:52]));

wire [5:0] layer1_N27_wire = {M0[323], M0[322], M0[309], M0[308], M0[65], M0[64]};
layer1_N27 layer1_N27_inst (.M0(layer1_N27_wire), .M1(M1[55:54]));

wire [5:0] layer1_N28_wire = {M0[471], M0[470], M0[257], M0[256], M0[145], M0[144]};
layer1_N28 layer1_N28_inst (.M0(layer1_N28_wire), .M1(M1[57:56]));

wire [5:0] layer1_N29_wire = {M0[259], M0[258], M0[221], M0[220], M0[75], M0[74]};
layer1_N29 layer1_N29_inst (.M0(layer1_N29_wire), .M1(M1[59:58]));

wire [5:0] layer1_N30_wire = {M0[347], M0[346], M0[321], M0[320], M0[47], M0[46]};
layer1_N30 layer1_N30_inst (.M0(layer1_N30_wire), .M1(M1[61:60]));

wire [5:0] layer1_N31_wire = {M0[479], M0[478], M0[311], M0[310], M0[67], M0[66]};
layer1_N31 layer1_N31_inst (.M0(layer1_N31_wire), .M1(M1[63:62]));

wire [5:0] layer1_N32_wire = {M0[405], M0[404], M0[345], M0[344], M0[9], M0[8]};
layer1_N32 layer1_N32_inst (.M0(layer1_N32_wire), .M1(M1[65:64]));

wire [5:0] layer1_N33_wire = {M0[505], M0[504], M0[481], M0[480], M0[141], M0[140]};
layer1_N33 layer1_N33_inst (.M0(layer1_N33_wire), .M1(M1[67:66]));

wire [5:0] layer1_N34_wire = {M0[411], M0[410], M0[329], M0[328], M0[131], M0[130]};
layer1_N34 layer1_N34_inst (.M0(layer1_N34_wire), .M1(M1[69:68]));

wire [5:0] layer1_N35_wire = {M0[421], M0[420], M0[219], M0[218], M0[61], M0[60]};
layer1_N35 layer1_N35_inst (.M0(layer1_N35_wire), .M1(M1[71:70]));

wire [5:0] layer1_N36_wire = {M0[487], M0[486], M0[483], M0[482], M0[163], M0[162]};
layer1_N36 layer1_N36_inst (.M0(layer1_N36_wire), .M1(M1[73:72]));

wire [5:0] layer1_N37_wire = {M0[309], M0[308], M0[277], M0[276], M0[31], M0[30]};
layer1_N37 layer1_N37_inst (.M0(layer1_N37_wire), .M1(M1[75:74]));

wire [5:0] layer1_N38_wire = {M0[343], M0[342], M0[317], M0[316], M0[21], M0[20]};
layer1_N38 layer1_N38_inst (.M0(layer1_N38_wire), .M1(M1[77:76]));

wire [5:0] layer1_N39_wire = {M0[481], M0[480], M0[385], M0[384], M0[259], M0[258]};
layer1_N39 layer1_N39_inst (.M0(layer1_N39_wire), .M1(M1[79:78]));

wire [5:0] layer1_N40_wire = {M0[465], M0[464], M0[243], M0[242], M0[45], M0[44]};
layer1_N40 layer1_N40_inst (.M0(layer1_N40_wire), .M1(M1[81:80]));

wire [5:0] layer1_N41_wire = {M0[335], M0[334], M0[305], M0[304], M0[241], M0[240]};
layer1_N41 layer1_N41_inst (.M0(layer1_N41_wire), .M1(M1[83:82]));

wire [5:0] layer1_N42_wire = {M0[223], M0[222], M0[219], M0[218], M0[181], M0[180]};
layer1_N42 layer1_N42_inst (.M0(layer1_N42_wire), .M1(M1[85:84]));

wire [5:0] layer1_N43_wire = {M0[461], M0[460], M0[281], M0[280], M0[101], M0[100]};
layer1_N43 layer1_N43_inst (.M0(layer1_N43_wire), .M1(M1[87:86]));

wire [5:0] layer1_N44_wire = {M0[459], M0[458], M0[349], M0[348], M0[271], M0[270]};
layer1_N44 layer1_N44_inst (.M0(layer1_N44_wire), .M1(M1[89:88]));

wire [5:0] layer1_N45_wire = {M0[209], M0[208], M0[41], M0[40], M0[37], M0[36]};
layer1_N45 layer1_N45_inst (.M0(layer1_N45_wire), .M1(M1[91:90]));

wire [5:0] layer1_N46_wire = {M0[423], M0[422], M0[369], M0[368], M0[157], M0[156]};
layer1_N46 layer1_N46_inst (.M0(layer1_N46_wire), .M1(M1[93:92]));

wire [5:0] layer1_N47_wire = {M0[343], M0[342], M0[213], M0[212], M0[31], M0[30]};
layer1_N47 layer1_N47_inst (.M0(layer1_N47_wire), .M1(M1[95:94]));

wire [5:0] layer1_N48_wire = {M0[305], M0[304], M0[121], M0[120], M0[87], M0[86]};
layer1_N48 layer1_N48_inst (.M0(layer1_N48_wire), .M1(M1[97:96]));

wire [5:0] layer1_N49_wire = {M0[391], M0[390], M0[163], M0[162], M0[121], M0[120]};
layer1_N49 layer1_N49_inst (.M0(layer1_N49_wire), .M1(M1[99:98]));

wire [5:0] layer1_N50_wire = {M0[413], M0[412], M0[313], M0[312], M0[253], M0[252]};
layer1_N50 layer1_N50_inst (.M0(layer1_N50_wire), .M1(M1[101:100]));

wire [5:0] layer1_N51_wire = {M0[363], M0[362], M0[251], M0[250], M0[53], M0[52]};
layer1_N51 layer1_N51_inst (.M0(layer1_N51_wire), .M1(M1[103:102]));

wire [5:0] layer1_N52_wire = {M0[469], M0[468], M0[331], M0[330], M0[217], M0[216]};
layer1_N52 layer1_N52_inst (.M0(layer1_N52_wire), .M1(M1[105:104]));

wire [5:0] layer1_N53_wire = {M0[411], M0[410], M0[305], M0[304], M0[297], M0[296]};
layer1_N53 layer1_N53_inst (.M0(layer1_N53_wire), .M1(M1[107:106]));

wire [5:0] layer1_N54_wire = {M0[429], M0[428], M0[213], M0[212], M0[57], M0[56]};
layer1_N54 layer1_N54_inst (.M0(layer1_N54_wire), .M1(M1[109:108]));

wire [5:0] layer1_N55_wire = {M0[427], M0[426], M0[179], M0[178], M0[63], M0[62]};
layer1_N55 layer1_N55_inst (.M0(layer1_N55_wire), .M1(M1[111:110]));

wire [5:0] layer1_N56_wire = {M0[207], M0[206], M0[89], M0[88], M0[31], M0[30]};
layer1_N56 layer1_N56_inst (.M0(layer1_N56_wire), .M1(M1[113:112]));

wire [5:0] layer1_N57_wire = {M0[485], M0[484], M0[443], M0[442], M0[141], M0[140]};
layer1_N57 layer1_N57_inst (.M0(layer1_N57_wire), .M1(M1[115:114]));

wire [5:0] layer1_N58_wire = {M0[449], M0[448], M0[47], M0[46], M0[1], M0[0]};
layer1_N58 layer1_N58_inst (.M0(layer1_N58_wire), .M1(M1[117:116]));

wire [5:0] layer1_N59_wire = {M0[503], M0[502], M0[455], M0[454], M0[251], M0[250]};
layer1_N59 layer1_N59_inst (.M0(layer1_N59_wire), .M1(M1[119:118]));

wire [5:0] layer1_N60_wire = {M0[479], M0[478], M0[303], M0[302], M0[117], M0[116]};
layer1_N60 layer1_N60_inst (.M0(layer1_N60_wire), .M1(M1[121:120]));

wire [5:0] layer1_N61_wire = {M0[389], M0[388], M0[341], M0[340], M0[187], M0[186]};
layer1_N61 layer1_N61_inst (.M0(layer1_N61_wire), .M1(M1[123:122]));

wire [5:0] layer1_N62_wire = {M0[153], M0[152], M0[125], M0[124], M0[23], M0[22]};
layer1_N62 layer1_N62_inst (.M0(layer1_N62_wire), .M1(M1[125:124]));

wire [5:0] layer1_N63_wire = {M0[489], M0[488], M0[209], M0[208], M0[39], M0[38]};
layer1_N63 layer1_N63_inst (.M0(layer1_N63_wire), .M1(M1[127:126]));

wire [5:0] layer1_N64_wire = {M0[461], M0[460], M0[285], M0[284], M0[275], M0[274]};
layer1_N64 layer1_N64_inst (.M0(layer1_N64_wire), .M1(M1[129:128]));

wire [5:0] layer1_N65_wire = {M0[511], M0[510], M0[399], M0[398], M0[29], M0[28]};
layer1_N65 layer1_N65_inst (.M0(layer1_N65_wire), .M1(M1[131:130]));

wire [5:0] layer1_N66_wire = {M0[435], M0[434], M0[187], M0[186], M0[33], M0[32]};
layer1_N66 layer1_N66_inst (.M0(layer1_N66_wire), .M1(M1[133:132]));

wire [5:0] layer1_N67_wire = {M0[313], M0[312], M0[117], M0[116], M0[99], M0[98]};
layer1_N67 layer1_N67_inst (.M0(layer1_N67_wire), .M1(M1[135:134]));

wire [5:0] layer1_N68_wire = {M0[171], M0[170], M0[125], M0[124], M0[115], M0[114]};
layer1_N68 layer1_N68_inst (.M0(layer1_N68_wire), .M1(M1[137:136]));

wire [5:0] layer1_N69_wire = {M0[225], M0[224], M0[175], M0[174], M0[153], M0[152]};
layer1_N69 layer1_N69_inst (.M0(layer1_N69_wire), .M1(M1[139:138]));

wire [5:0] layer1_N70_wire = {M0[361], M0[360], M0[327], M0[326], M0[103], M0[102]};
layer1_N70 layer1_N70_inst (.M0(layer1_N70_wire), .M1(M1[141:140]));

wire [5:0] layer1_N71_wire = {M0[91], M0[90], M0[37], M0[36], M0[25], M0[24]};
layer1_N71 layer1_N71_inst (.M0(layer1_N71_wire), .M1(M1[143:142]));

wire [5:0] layer1_N72_wire = {M0[453], M0[452], M0[247], M0[246], M0[93], M0[92]};
layer1_N72 layer1_N72_inst (.M0(layer1_N72_wire), .M1(M1[145:144]));

wire [5:0] layer1_N73_wire = {M0[511], M0[510], M0[481], M0[480], M0[295], M0[294]};
layer1_N73 layer1_N73_inst (.M0(layer1_N73_wire), .M1(M1[147:146]));

wire [5:0] layer1_N74_wire = {M0[347], M0[346], M0[329], M0[328], M0[305], M0[304]};
layer1_N74 layer1_N74_inst (.M0(layer1_N74_wire), .M1(M1[149:148]));

wire [5:0] layer1_N75_wire = {M0[89], M0[88], M0[63], M0[62], M0[47], M0[46]};
layer1_N75 layer1_N75_inst (.M0(layer1_N75_wire), .M1(M1[151:150]));

wire [5:0] layer1_N76_wire = {M0[459], M0[458], M0[247], M0[246], M0[7], M0[6]};
layer1_N76 layer1_N76_inst (.M0(layer1_N76_wire), .M1(M1[153:152]));

wire [5:0] layer1_N77_wire = {M0[453], M0[452], M0[445], M0[444], M0[61], M0[60]};
layer1_N77 layer1_N77_inst (.M0(layer1_N77_wire), .M1(M1[155:154]));

wire [5:0] layer1_N78_wire = {M0[329], M0[328], M0[203], M0[202], M0[149], M0[148]};
layer1_N78 layer1_N78_inst (.M0(layer1_N78_wire), .M1(M1[157:156]));

wire [5:0] layer1_N79_wire = {M0[369], M0[368], M0[343], M0[342], M0[237], M0[236]};
layer1_N79 layer1_N79_inst (.M0(layer1_N79_wire), .M1(M1[159:158]));

wire [5:0] layer1_N80_wire = {M0[249], M0[248], M0[205], M0[204], M0[153], M0[152]};
layer1_N80 layer1_N80_inst (.M0(layer1_N80_wire), .M1(M1[161:160]));

wire [5:0] layer1_N81_wire = {M0[349], M0[348], M0[117], M0[116], M0[39], M0[38]};
layer1_N81 layer1_N81_inst (.M0(layer1_N81_wire), .M1(M1[163:162]));

wire [5:0] layer1_N82_wire = {M0[475], M0[474], M0[149], M0[148], M0[31], M0[30]};
layer1_N82 layer1_N82_inst (.M0(layer1_N82_wire), .M1(M1[165:164]));

wire [5:0] layer1_N83_wire = {M0[155], M0[154], M0[105], M0[104], M0[35], M0[34]};
layer1_N83 layer1_N83_inst (.M0(layer1_N83_wire), .M1(M1[167:166]));

wire [5:0] layer1_N84_wire = {M0[511], M0[510], M0[253], M0[252], M0[119], M0[118]};
layer1_N84 layer1_N84_inst (.M0(layer1_N84_wire), .M1(M1[169:168]));

wire [5:0] layer1_N85_wire = {M0[259], M0[258], M0[95], M0[94], M0[93], M0[92]};
layer1_N85 layer1_N85_inst (.M0(layer1_N85_wire), .M1(M1[171:170]));

endmodule