module layer0 (input [511:0] M0, output [511:0] M1);

wire [5:0] layer0_N0_wire = {M0[474], M0[384], M0[353], M0[262], M0[40], M0[27]};
layer0_N0 layer0_N0_inst (.M0(layer0_N0_wire), .M1(M1[1:0]));

wire [5:0] layer0_N1_wire = {M0[436], M0[398], M0[270], M0[161], M0[74], M0[48]};
layer0_N1 layer0_N1_inst (.M0(layer0_N1_wire), .M1(M1[3:2]));

wire [5:0] layer0_N2_wire = {M0[467], M0[435], M0[421], M0[163], M0[143], M0[95]};
layer0_N2 layer0_N2_inst (.M0(layer0_N2_wire), .M1(M1[5:4]));

wire [5:0] layer0_N3_wire = {M0[500], M0[382], M0[315], M0[284], M0[220], M0[37]};
layer0_N3 layer0_N3_inst (.M0(layer0_N3_wire), .M1(M1[7:6]));

wire [5:0] layer0_N4_wire = {M0[404], M0[299], M0[79], M0[33], M0[20], M0[4]};
layer0_N4 layer0_N4_inst (.M0(layer0_N4_wire), .M1(M1[9:8]));

wire [5:0] layer0_N5_wire = {M0[509], M0[441], M0[388], M0[254], M0[66], M0[48]};
layer0_N5 layer0_N5_inst (.M0(layer0_N5_wire), .M1(M1[11:10]));

wire [5:0] layer0_N6_wire = {M0[497], M0[494], M0[249], M0[239], M0[194], M0[64]};
layer0_N6 layer0_N6_inst (.M0(layer0_N6_wire), .M1(M1[13:12]));

wire [5:0] layer0_N7_wire = {M0[461], M0[412], M0[356], M0[164], M0[142], M0[100]};
layer0_N7 layer0_N7_inst (.M0(layer0_N7_wire), .M1(M1[15:14]));

wire [5:0] layer0_N8_wire = {M0[457], M0[403], M0[382], M0[225], M0[89], M0[61]};
layer0_N8 layer0_N8_inst (.M0(layer0_N8_wire), .M1(M1[17:16]));

wire [5:0] layer0_N9_wire = {M0[490], M0[472], M0[400], M0[375], M0[103], M0[14]};
layer0_N9 layer0_N9_inst (.M0(layer0_N9_wire), .M1(M1[19:18]));

wire [5:0] layer0_N10_wire = {M0[486], M0[410], M0[359], M0[48], M0[32], M0[31]};
layer0_N10 layer0_N10_inst (.M0(layer0_N10_wire), .M1(M1[21:20]));

wire [5:0] layer0_N11_wire = {M0[433], M0[372], M0[262], M0[225], M0[151], M0[13]};
layer0_N11 layer0_N11_inst (.M0(layer0_N11_wire), .M1(M1[23:22]));

wire [5:0] layer0_N12_wire = {M0[474], M0[452], M0[343], M0[284], M0[89], M0[13]};
layer0_N12 layer0_N12_inst (.M0(layer0_N12_wire), .M1(M1[25:24]));

wire [5:0] layer0_N13_wire = {M0[427], M0[328], M0[322], M0[227], M0[197], M0[136]};
layer0_N13 layer0_N13_inst (.M0(layer0_N13_wire), .M1(M1[27:26]));

wire [5:0] layer0_N14_wire = {M0[503], M0[348], M0[274], M0[161], M0[154], M0[152]};
layer0_N14 layer0_N14_inst (.M0(layer0_N14_wire), .M1(M1[29:28]));

wire [5:0] layer0_N15_wire = {M0[477], M0[474], M0[440], M0[409], M0[395], M0[152]};
layer0_N15 layer0_N15_inst (.M0(layer0_N15_wire), .M1(M1[31:30]));

wire [5:0] layer0_N16_wire = {M0[403], M0[389], M0[388], M0[381], M0[268], M0[201]};
layer0_N16 layer0_N16_inst (.M0(layer0_N16_wire), .M1(M1[33:32]));

wire [5:0] layer0_N17_wire = {M0[486], M0[424], M0[346], M0[268], M0[168], M0[150]};
layer0_N17 layer0_N17_inst (.M0(layer0_N17_wire), .M1(M1[35:34]));

wire [5:0] layer0_N18_wire = {M0[391], M0[375], M0[266], M0[197], M0[40], M0[7]};
layer0_N18 layer0_N18_inst (.M0(layer0_N18_wire), .M1(M1[37:36]));

wire [5:0] layer0_N19_wire = {M0[506], M0[434], M0[318], M0[247], M0[191], M0[176]};
layer0_N19 layer0_N19_inst (.M0(layer0_N19_wire), .M1(M1[39:38]));

wire [5:0] layer0_N20_wire = {M0[463], M0[278], M0[243], M0[206], M0[154], M0[147]};
layer0_N20 layer0_N20_inst (.M0(layer0_N20_wire), .M1(M1[41:40]));

wire [5:0] layer0_N21_wire = {M0[456], M0[452], M0[196], M0[168], M0[95], M0[54]};
layer0_N21 layer0_N21_inst (.M0(layer0_N21_wire), .M1(M1[43:42]));

wire [5:0] layer0_N22_wire = {M0[472], M0[350], M0[281], M0[237], M0[230], M0[6]};
layer0_N22 layer0_N22_inst (.M0(layer0_N22_wire), .M1(M1[45:44]));

wire [5:0] layer0_N23_wire = {M0[408], M0[189], M0[146], M0[137], M0[81], M0[80]};
layer0_N23 layer0_N23_inst (.M0(layer0_N23_wire), .M1(M1[47:46]));

wire [5:0] layer0_N24_wire = {M0[455], M0[440], M0[415], M0[412], M0[342], M0[147]};
layer0_N24 layer0_N24_inst (.M0(layer0_N24_wire), .M1(M1[49:48]));

wire [5:0] layer0_N25_wire = {M0[473], M0[451], M0[446], M0[333], M0[172], M0[48]};
layer0_N25 layer0_N25_inst (.M0(layer0_N25_wire), .M1(M1[51:50]));

wire [5:0] layer0_N26_wire = {M0[508], M0[505], M0[212], M0[172], M0[158], M0[5]};
layer0_N26 layer0_N26_inst (.M0(layer0_N26_wire), .M1(M1[53:52]));

wire [5:0] layer0_N27_wire = {M0[245], M0[225], M0[157], M0[113], M0[68], M0[47]};
layer0_N27 layer0_N27_inst (.M0(layer0_N27_wire), .M1(M1[55:54]));

wire [5:0] layer0_N28_wire = {M0[361], M0[345], M0[316], M0[269], M0[168], M0[129]};
layer0_N28 layer0_N28_inst (.M0(layer0_N28_wire), .M1(M1[57:56]));

wire [5:0] layer0_N29_wire = {M0[490], M0[275], M0[196], M0[117], M0[95], M0[39]};
layer0_N29 layer0_N29_inst (.M0(layer0_N29_wire), .M1(M1[59:58]));

wire [5:0] layer0_N30_wire = {M0[500], M0[486], M0[450], M0[418], M0[172], M0[75]};
layer0_N30 layer0_N30_inst (.M0(layer0_N30_wire), .M1(M1[61:60]));

wire [5:0] layer0_N31_wire = {M0[510], M0[435], M0[328], M0[323], M0[267], M0[52]};
layer0_N31 layer0_N31_inst (.M0(layer0_N31_wire), .M1(M1[63:62]));

wire [5:0] layer0_N32_wire = {M0[270], M0[242], M0[179], M0[66], M0[61], M0[26]};
layer0_N32 layer0_N32_inst (.M0(layer0_N32_wire), .M1(M1[65:64]));

wire [5:0] layer0_N33_wire = {M0[467], M0[445], M0[425], M0[225], M0[170], M0[134]};
layer0_N33 layer0_N33_inst (.M0(layer0_N33_wire), .M1(M1[67:66]));

wire [5:0] layer0_N34_wire = {M0[494], M0[402], M0[308], M0[289], M0[198], M0[195]};
layer0_N34 layer0_N34_inst (.M0(layer0_N34_wire), .M1(M1[69:68]));

wire [5:0] layer0_N35_wire = {M0[503], M0[336], M0[254], M0[78], M0[57], M0[53]};
layer0_N35 layer0_N35_inst (.M0(layer0_N35_wire), .M1(M1[71:70]));

wire [5:0] layer0_N36_wire = {M0[500], M0[457], M0[372], M0[306], M0[257], M0[81]};
layer0_N36 layer0_N36_inst (.M0(layer0_N36_wire), .M1(M1[73:72]));

wire [5:0] layer0_N37_wire = {M0[416], M0[339], M0[156], M0[108], M0[81], M0[40]};
layer0_N37 layer0_N37_inst (.M0(layer0_N37_wire), .M1(M1[75:74]));

wire [5:0] layer0_N38_wire = {M0[429], M0[402], M0[259], M0[206], M0[130], M0[39]};
layer0_N38 layer0_N38_inst (.M0(layer0_N38_wire), .M1(M1[77:76]));

wire [5:0] layer0_N39_wire = {M0[507], M0[500], M0[452], M0[263], M0[36], M0[32]};
layer0_N39 layer0_N39_inst (.M0(layer0_N39_wire), .M1(M1[79:78]));

wire [5:0] layer0_N40_wire = {M0[403], M0[350], M0[332], M0[223], M0[216], M0[0]};
layer0_N40 layer0_N40_inst (.M0(layer0_N40_wire), .M1(M1[81:80]));

wire [5:0] layer0_N41_wire = {M0[511], M0[326], M0[176], M0[72], M0[64], M0[20]};
layer0_N41 layer0_N41_inst (.M0(layer0_N41_wire), .M1(M1[83:82]));

wire [5:0] layer0_N42_wire = {M0[437], M0[395], M0[337], M0[307], M0[93], M0[87]};
layer0_N42 layer0_N42_inst (.M0(layer0_N42_wire), .M1(M1[85:84]));

wire [5:0] layer0_N43_wire = {M0[495], M0[493], M0[306], M0[182], M0[157], M0[33]};
layer0_N43 layer0_N43_inst (.M0(layer0_N43_wire), .M1(M1[87:86]));

wire [5:0] layer0_N44_wire = {M0[509], M0[371], M0[257], M0[164], M0[121], M0[16]};
layer0_N44 layer0_N44_inst (.M0(layer0_N44_wire), .M1(M1[89:88]));

wire [5:0] layer0_N45_wire = {M0[337], M0[207], M0[183], M0[94], M0[63], M0[32]};
layer0_N45 layer0_N45_inst (.M0(layer0_N45_wire), .M1(M1[91:90]));

wire [5:0] layer0_N46_wire = {M0[323], M0[306], M0[301], M0[159], M0[139], M0[39]};
layer0_N46 layer0_N46_inst (.M0(layer0_N46_wire), .M1(M1[93:92]));

wire [5:0] layer0_N47_wire = {M0[490], M0[427], M0[122], M0[71], M0[61], M0[34]};
layer0_N47 layer0_N47_inst (.M0(layer0_N47_wire), .M1(M1[95:94]));

wire [5:0] layer0_N48_wire = {M0[457], M0[437], M0[398], M0[255], M0[248], M0[99]};
layer0_N48 layer0_N48_inst (.M0(layer0_N48_wire), .M1(M1[97:96]));

wire [5:0] layer0_N49_wire = {M0[459], M0[362], M0[234], M0[223], M0[171], M0[54]};
layer0_N49 layer0_N49_inst (.M0(layer0_N49_wire), .M1(M1[99:98]));

wire [5:0] layer0_N50_wire = {M0[296], M0[271], M0[270], M0[263], M0[21], M0[18]};
layer0_N50 layer0_N50_inst (.M0(layer0_N50_wire), .M1(M1[101:100]));

wire [5:0] layer0_N51_wire = {M0[483], M0[479], M0[304], M0[138], M0[131], M0[82]};
layer0_N51 layer0_N51_inst (.M0(layer0_N51_wire), .M1(M1[103:102]));

wire [5:0] layer0_N52_wire = {M0[511], M0[456], M0[240], M0[208], M0[126], M0[90]};
layer0_N52 layer0_N52_inst (.M0(layer0_N52_wire), .M1(M1[105:104]));

wire [5:0] layer0_N53_wire = {M0[433], M0[344], M0[239], M0[169], M0[161], M0[99]};
layer0_N53 layer0_N53_inst (.M0(layer0_N53_wire), .M1(M1[107:106]));

wire [5:0] layer0_N54_wire = {M0[476], M0[352], M0[242], M0[98], M0[33], M0[9]};
layer0_N54 layer0_N54_inst (.M0(layer0_N54_wire), .M1(M1[109:108]));

wire [5:0] layer0_N55_wire = {M0[500], M0[328], M0[282], M0[102], M0[61], M0[57]};
layer0_N55 layer0_N55_inst (.M0(layer0_N55_wire), .M1(M1[111:110]));

wire [5:0] layer0_N56_wire = {M0[406], M0[384], M0[294], M0[77], M0[67], M0[11]};
layer0_N56 layer0_N56_inst (.M0(layer0_N56_wire), .M1(M1[113:112]));

wire [5:0] layer0_N57_wire = {M0[421], M0[407], M0[328], M0[296], M0[275], M0[163]};
layer0_N57 layer0_N57_inst (.M0(layer0_N57_wire), .M1(M1[115:114]));

wire [5:0] layer0_N58_wire = {M0[488], M0[475], M0[441], M0[397], M0[331], M0[100]};
layer0_N58 layer0_N58_inst (.M0(layer0_N58_wire), .M1(M1[117:116]));

wire [5:0] layer0_N59_wire = {M0[444], M0[424], M0[348], M0[190], M0[170], M0[167]};
layer0_N59 layer0_N59_inst (.M0(layer0_N59_wire), .M1(M1[119:118]));

wire [5:0] layer0_N60_wire = {M0[504], M0[495], M0[472], M0[288], M0[138], M0[82]};
layer0_N60 layer0_N60_inst (.M0(layer0_N60_wire), .M1(M1[121:120]));

wire [5:0] layer0_N61_wire = {M0[393], M0[232], M0[198], M0[167], M0[58], M0[3]};
layer0_N61 layer0_N61_inst (.M0(layer0_N61_wire), .M1(M1[123:122]));

wire [5:0] layer0_N62_wire = {M0[472], M0[424], M0[418], M0[383], M0[351], M0[99]};
layer0_N62 layer0_N62_inst (.M0(layer0_N62_wire), .M1(M1[125:124]));

wire [5:0] layer0_N63_wire = {M0[447], M0[407], M0[227], M0[150], M0[124], M0[55]};
layer0_N63 layer0_N63_inst (.M0(layer0_N63_wire), .M1(M1[127:126]));

wire [5:0] layer0_N64_wire = {M0[438], M0[370], M0[288], M0[283], M0[226], M0[37]};
layer0_N64 layer0_N64_inst (.M0(layer0_N64_wire), .M1(M1[129:128]));

wire [5:0] layer0_N65_wire = {M0[441], M0[317], M0[248], M0[202], M0[93], M0[80]};
layer0_N65 layer0_N65_inst (.M0(layer0_N65_wire), .M1(M1[131:130]));

wire [5:0] layer0_N66_wire = {M0[457], M0[277], M0[273], M0[250], M0[234], M0[49]};
layer0_N66 layer0_N66_inst (.M0(layer0_N66_wire), .M1(M1[133:132]));

wire [5:0] layer0_N67_wire = {M0[492], M0[443], M0[442], M0[402], M0[208], M0[38]};
layer0_N67 layer0_N67_inst (.M0(layer0_N67_wire), .M1(M1[135:134]));

wire [5:0] layer0_N68_wire = {M0[428], M0[409], M0[279], M0[247], M0[179], M0[43]};
layer0_N68 layer0_N68_inst (.M0(layer0_N68_wire), .M1(M1[137:136]));

wire [5:0] layer0_N69_wire = {M0[449], M0[390], M0[306], M0[96], M0[83], M0[24]};
layer0_N69 layer0_N69_inst (.M0(layer0_N69_wire), .M1(M1[139:138]));

wire [5:0] layer0_N70_wire = {M0[500], M0[457], M0[218], M0[146], M0[134], M0[47]};
layer0_N70 layer0_N70_inst (.M0(layer0_N70_wire), .M1(M1[141:140]));

wire [5:0] layer0_N71_wire = {M0[511], M0[355], M0[264], M0[216], M0[211], M0[201]};
layer0_N71 layer0_N71_inst (.M0(layer0_N71_wire), .M1(M1[143:142]));

wire [5:0] layer0_N72_wire = {M0[486], M0[416], M0[209], M0[91], M0[65], M0[52]};
layer0_N72 layer0_N72_inst (.M0(layer0_N72_wire), .M1(M1[145:144]));

wire [5:0] layer0_N73_wire = {M0[491], M0[345], M0[259], M0[194], M0[178], M0[32]};
layer0_N73 layer0_N73_inst (.M0(layer0_N73_wire), .M1(M1[147:146]));

wire [5:0] layer0_N74_wire = {M0[504], M0[469], M0[327], M0[312], M0[293], M0[49]};
layer0_N74 layer0_N74_inst (.M0(layer0_N74_wire), .M1(M1[149:148]));

wire [5:0] layer0_N75_wire = {M0[422], M0[258], M0[93], M0[72], M0[70], M0[24]};
layer0_N75 layer0_N75_inst (.M0(layer0_N75_wire), .M1(M1[151:150]));

wire [5:0] layer0_N76_wire = {M0[381], M0[375], M0[350], M0[347], M0[157], M0[122]};
layer0_N76 layer0_N76_inst (.M0(layer0_N76_wire), .M1(M1[153:152]));

wire [5:0] layer0_N77_wire = {M0[425], M0[363], M0[334], M0[298], M0[202], M0[161]};
layer0_N77 layer0_N77_inst (.M0(layer0_N77_wire), .M1(M1[155:154]));

wire [5:0] layer0_N78_wire = {M0[257], M0[234], M0[176], M0[42], M0[33], M0[21]};
layer0_N78 layer0_N78_inst (.M0(layer0_N78_wire), .M1(M1[157:156]));

wire [5:0] layer0_N79_wire = {M0[234], M0[224], M0[156], M0[119], M0[90], M0[26]};
layer0_N79 layer0_N79_inst (.M0(layer0_N79_wire), .M1(M1[159:158]));

wire [5:0] layer0_N80_wire = {M0[482], M0[476], M0[448], M0[371], M0[233], M0[62]};
layer0_N80 layer0_N80_inst (.M0(layer0_N80_wire), .M1(M1[161:160]));

wire [5:0] layer0_N81_wire = {M0[456], M0[451], M0[392], M0[379], M0[98], M0[38]};
layer0_N81 layer0_N81_inst (.M0(layer0_N81_wire), .M1(M1[163:162]));

wire [5:0] layer0_N82_wire = {M0[470], M0[420], M0[166], M0[157], M0[144], M0[8]};
layer0_N82 layer0_N82_inst (.M0(layer0_N82_wire), .M1(M1[165:164]));

wire [5:0] layer0_N83_wire = {M0[468], M0[341], M0[274], M0[217], M0[152], M0[52]};
layer0_N83 layer0_N83_inst (.M0(layer0_N83_wire), .M1(M1[167:166]));

wire [5:0] layer0_N84_wire = {M0[399], M0[252], M0[247], M0[236], M0[116], M0[64]};
layer0_N84 layer0_N84_inst (.M0(layer0_N84_wire), .M1(M1[169:168]));

wire [5:0] layer0_N85_wire = {M0[382], M0[365], M0[324], M0[81], M0[51], M0[26]};
layer0_N85 layer0_N85_inst (.M0(layer0_N85_wire), .M1(M1[171:170]));

wire [5:0] layer0_N86_wire = {M0[501], M0[368], M0[343], M0[213], M0[82], M0[53]};
layer0_N86 layer0_N86_inst (.M0(layer0_N86_wire), .M1(M1[173:172]));

wire [5:0] layer0_N87_wire = {M0[480], M0[435], M0[384], M0[314], M0[285], M0[24]};
layer0_N87 layer0_N87_inst (.M0(layer0_N87_wire), .M1(M1[175:174]));

wire [5:0] layer0_N88_wire = {M0[450], M0[420], M0[290], M0[270], M0[90], M0[54]};
layer0_N88 layer0_N88_inst (.M0(layer0_N88_wire), .M1(M1[177:176]));

wire [5:0] layer0_N89_wire = {M0[496], M0[436], M0[412], M0[305], M0[228], M0[134]};
layer0_N89 layer0_N89_inst (.M0(layer0_N89_wire), .M1(M1[179:178]));

wire [5:0] layer0_N90_wire = {M0[505], M0[453], M0[446], M0[197], M0[158], M0[148]};
layer0_N90 layer0_N90_inst (.M0(layer0_N90_wire), .M1(M1[181:180]));

wire [5:0] layer0_N91_wire = {M0[462], M0[436], M0[345], M0[340], M0[319], M0[56]};
layer0_N91 layer0_N91_inst (.M0(layer0_N91_wire), .M1(M1[183:182]));

wire [5:0] layer0_N92_wire = {M0[407], M0[237], M0[186], M0[141], M0[77], M0[0]};
layer0_N92 layer0_N92_inst (.M0(layer0_N92_wire), .M1(M1[185:184]));

wire [5:0] layer0_N93_wire = {M0[436], M0[257], M0[224], M0[216], M0[173], M0[97]};
layer0_N93 layer0_N93_inst (.M0(layer0_N93_wire), .M1(M1[187:186]));

wire [5:0] layer0_N94_wire = {M0[484], M0[477], M0[443], M0[397], M0[344], M0[13]};
layer0_N94 layer0_N94_inst (.M0(layer0_N94_wire), .M1(M1[189:188]));

wire [5:0] layer0_N95_wire = {M0[284], M0[224], M0[150], M0[146], M0[138], M0[54]};
layer0_N95 layer0_N95_inst (.M0(layer0_N95_wire), .M1(M1[191:190]));

wire [5:0] layer0_N96_wire = {M0[221], M0[161], M0[120], M0[68], M0[44], M0[16]};
layer0_N96 layer0_N96_inst (.M0(layer0_N96_wire), .M1(M1[193:192]));

wire [5:0] layer0_N97_wire = {M0[469], M0[368], M0[283], M0[273], M0[247], M0[85]};
layer0_N97 layer0_N97_inst (.M0(layer0_N97_wire), .M1(M1[195:194]));

wire [5:0] layer0_N98_wire = {M0[432], M0[404], M0[201], M0[118], M0[35], M0[24]};
layer0_N98 layer0_N98_inst (.M0(layer0_N98_wire), .M1(M1[197:196]));

wire [5:0] layer0_N99_wire = {M0[510], M0[335], M0[157], M0[155], M0[64], M0[16]};
layer0_N99 layer0_N99_inst (.M0(layer0_N99_wire), .M1(M1[199:198]));

wire [5:0] layer0_N100_wire = {M0[467], M0[417], M0[305], M0[289], M0[110], M0[62]};
layer0_N100 layer0_N100_inst (.M0(layer0_N100_wire), .M1(M1[201:200]));

wire [5:0] layer0_N101_wire = {M0[440], M0[385], M0[276], M0[144], M0[125], M0[17]};
layer0_N101 layer0_N101_inst (.M0(layer0_N101_wire), .M1(M1[203:202]));

wire [5:0] layer0_N102_wire = {M0[377], M0[369], M0[302], M0[237], M0[53], M0[9]};
layer0_N102 layer0_N102_inst (.M0(layer0_N102_wire), .M1(M1[205:204]));

wire [5:0] layer0_N103_wire = {M0[511], M0[460], M0[357], M0[329], M0[150], M0[19]};
layer0_N103 layer0_N103_inst (.M0(layer0_N103_wire), .M1(M1[207:206]));

wire [5:0] layer0_N104_wire = {M0[407], M0[341], M0[237], M0[207], M0[112], M0[77]};
layer0_N104 layer0_N104_inst (.M0(layer0_N104_wire), .M1(M1[209:208]));

wire [5:0] layer0_N105_wire = {M0[334], M0[318], M0[289], M0[286], M0[208], M0[192]};
layer0_N105 layer0_N105_inst (.M0(layer0_N105_wire), .M1(M1[211:210]));

wire [5:0] layer0_N106_wire = {M0[490], M0[464], M0[446], M0[438], M0[296], M0[187]};
layer0_N106 layer0_N106_inst (.M0(layer0_N106_wire), .M1(M1[213:212]));

wire [5:0] layer0_N107_wire = {M0[433], M0[320], M0[304], M0[273], M0[162], M0[150]};
layer0_N107 layer0_N107_inst (.M0(layer0_N107_wire), .M1(M1[215:214]));

wire [5:0] layer0_N108_wire = {M0[452], M0[419], M0[391], M0[373], M0[142], M0[33]};
layer0_N108 layer0_N108_inst (.M0(layer0_N108_wire), .M1(M1[217:216]));

wire [5:0] layer0_N109_wire = {M0[470], M0[422], M0[410], M0[356], M0[150], M0[85]};
layer0_N109 layer0_N109_inst (.M0(layer0_N109_wire), .M1(M1[219:218]));

wire [5:0] layer0_N110_wire = {M0[507], M0[321], M0[281], M0[218], M0[216], M0[71]};
layer0_N110 layer0_N110_inst (.M0(layer0_N110_wire), .M1(M1[221:220]));

wire [5:0] layer0_N111_wire = {M0[509], M0[488], M0[383], M0[208], M0[148], M0[2]};
layer0_N111 layer0_N111_inst (.M0(layer0_N111_wire), .M1(M1[223:222]));

wire [5:0] layer0_N112_wire = {M0[435], M0[380], M0[217], M0[130], M0[68], M0[35]};
layer0_N112 layer0_N112_inst (.M0(layer0_N112_wire), .M1(M1[225:224]));

wire [5:0] layer0_N113_wire = {M0[484], M0[469], M0[113], M0[101], M0[83], M0[4]};
layer0_N113 layer0_N113_inst (.M0(layer0_N113_wire), .M1(M1[227:226]));

wire [5:0] layer0_N114_wire = {M0[379], M0[329], M0[310], M0[302], M0[149], M0[89]};
layer0_N114 layer0_N114_inst (.M0(layer0_N114_wire), .M1(M1[229:228]));

wire [5:0] layer0_N115_wire = {M0[399], M0[356], M0[351], M0[348], M0[318], M0[98]};
layer0_N115 layer0_N115_inst (.M0(layer0_N115_wire), .M1(M1[231:230]));

wire [5:0] layer0_N116_wire = {M0[499], M0[403], M0[292], M0[279], M0[187], M0[182]};
layer0_N116 layer0_N116_inst (.M0(layer0_N116_wire), .M1(M1[233:232]));

wire [5:0] layer0_N117_wire = {M0[504], M0[351], M0[343], M0[222], M0[206], M0[79]};
layer0_N117 layer0_N117_inst (.M0(layer0_N117_wire), .M1(M1[235:234]));

wire [5:0] layer0_N118_wire = {M0[393], M0[240], M0[205], M0[72], M0[55], M0[7]};
layer0_N118 layer0_N118_inst (.M0(layer0_N118_wire), .M1(M1[237:236]));

wire [5:0] layer0_N119_wire = {M0[489], M0[354], M0[177], M0[95], M0[81], M0[71]};
layer0_N119 layer0_N119_inst (.M0(layer0_N119_wire), .M1(M1[239:238]));

wire [5:0] layer0_N120_wire = {M0[484], M0[461], M0[160], M0[73], M0[57], M0[16]};
layer0_N120 layer0_N120_inst (.M0(layer0_N120_wire), .M1(M1[241:240]));

wire [5:0] layer0_N121_wire = {M0[446], M0[413], M0[324], M0[311], M0[286], M0[2]};
layer0_N121 layer0_N121_inst (.M0(layer0_N121_wire), .M1(M1[243:242]));

wire [5:0] layer0_N122_wire = {M0[413], M0[284], M0[260], M0[258], M0[119], M0[49]};
layer0_N122 layer0_N122_inst (.M0(layer0_N122_wire), .M1(M1[245:244]));

wire [5:0] layer0_N123_wire = {M0[444], M0[314], M0[298], M0[237], M0[216], M0[29]};
layer0_N123 layer0_N123_inst (.M0(layer0_N123_wire), .M1(M1[247:246]));

wire [5:0] layer0_N124_wire = {M0[438], M0[404], M0[392], M0[372], M0[245], M0[194]};
layer0_N124 layer0_N124_inst (.M0(layer0_N124_wire), .M1(M1[249:248]));

wire [5:0] layer0_N125_wire = {M0[463], M0[392], M0[177], M0[97], M0[43], M0[21]};
layer0_N125 layer0_N125_inst (.M0(layer0_N125_wire), .M1(M1[251:250]));

wire [5:0] layer0_N126_wire = {M0[462], M0[461], M0[347], M0[322], M0[302], M0[223]};
layer0_N126 layer0_N126_inst (.M0(layer0_N126_wire), .M1(M1[253:252]));

wire [5:0] layer0_N127_wire = {M0[444], M0[386], M0[336], M0[245], M0[228], M0[15]};
layer0_N127 layer0_N127_inst (.M0(layer0_N127_wire), .M1(M1[255:254]));

wire [5:0] layer0_N128_wire = {M0[341], M0[301], M0[259], M0[249], M0[238], M0[112]};
layer0_N128 layer0_N128_inst (.M0(layer0_N128_wire), .M1(M1[257:256]));

wire [5:0] layer0_N129_wire = {M0[360], M0[336], M0[327], M0[127], M0[82], M0[76]};
layer0_N129 layer0_N129_inst (.M0(layer0_N129_wire), .M1(M1[259:258]));

wire [5:0] layer0_N130_wire = {M0[500], M0[358], M0[283], M0[270], M0[51], M0[46]};
layer0_N130 layer0_N130_inst (.M0(layer0_N130_wire), .M1(M1[261:260]));

wire [5:0] layer0_N131_wire = {M0[501], M0[483], M0[342], M0[285], M0[231], M0[201]};
layer0_N131 layer0_N131_inst (.M0(layer0_N131_wire), .M1(M1[263:262]));

wire [5:0] layer0_N132_wire = {M0[400], M0[360], M0[343], M0[295], M0[165], M0[90]};
layer0_N132 layer0_N132_inst (.M0(layer0_N132_wire), .M1(M1[265:264]));

wire [5:0] layer0_N133_wire = {M0[385], M0[372], M0[287], M0[246], M0[174], M0[59]};
layer0_N133 layer0_N133_inst (.M0(layer0_N133_wire), .M1(M1[267:266]));

wire [5:0] layer0_N134_wire = {M0[300], M0[252], M0[171], M0[82], M0[69], M0[64]};
layer0_N134 layer0_N134_inst (.M0(layer0_N134_wire), .M1(M1[269:268]));

wire [5:0] layer0_N135_wire = {M0[511], M0[488], M0[269], M0[248], M0[239], M0[36]};
layer0_N135 layer0_N135_inst (.M0(layer0_N135_wire), .M1(M1[271:270]));

wire [5:0] layer0_N136_wire = {M0[398], M0[325], M0[257], M0[188], M0[128], M0[44]};
layer0_N136 layer0_N136_inst (.M0(layer0_N136_wire), .M1(M1[273:272]));

wire [5:0] layer0_N137_wire = {M0[457], M0[311], M0[308], M0[221], M0[168], M0[94]};
layer0_N137 layer0_N137_inst (.M0(layer0_N137_wire), .M1(M1[275:274]));

wire [5:0] layer0_N138_wire = {M0[500], M0[397], M0[319], M0[307], M0[139], M0[83]};
layer0_N138 layer0_N138_inst (.M0(layer0_N138_wire), .M1(M1[277:276]));

wire [5:0] layer0_N139_wire = {M0[480], M0[473], M0[268], M0[238], M0[219], M0[70]};
layer0_N139 layer0_N139_inst (.M0(layer0_N139_wire), .M1(M1[279:278]));

wire [5:0] layer0_N140_wire = {M0[490], M0[353], M0[299], M0[201], M0[183], M0[133]};
layer0_N140 layer0_N140_inst (.M0(layer0_N140_wire), .M1(M1[281:280]));

wire [5:0] layer0_N141_wire = {M0[492], M0[419], M0[353], M0[103], M0[32], M0[10]};
layer0_N141 layer0_N141_inst (.M0(layer0_N141_wire), .M1(M1[283:282]));

wire [5:0] layer0_N142_wire = {M0[432], M0[389], M0[354], M0[236], M0[111], M0[26]};
layer0_N142 layer0_N142_inst (.M0(layer0_N142_wire), .M1(M1[285:284]));

wire [5:0] layer0_N143_wire = {M0[470], M0[285], M0[258], M0[228], M0[41], M0[40]};
layer0_N143 layer0_N143_inst (.M0(layer0_N143_wire), .M1(M1[287:286]));

wire [5:0] layer0_N144_wire = {M0[487], M0[452], M0[427], M0[404], M0[329], M0[50]};
layer0_N144 layer0_N144_inst (.M0(layer0_N144_wire), .M1(M1[289:288]));

wire [5:0] layer0_N145_wire = {M0[425], M0[301], M0[168], M0[152], M0[130], M0[126]};
layer0_N145 layer0_N145_inst (.M0(layer0_N145_wire), .M1(M1[291:290]));

wire [5:0] layer0_N146_wire = {M0[440], M0[223], M0[208], M0[200], M0[195], M0[15]};
layer0_N146 layer0_N146_inst (.M0(layer0_N146_wire), .M1(M1[293:292]));

wire [5:0] layer0_N147_wire = {M0[462], M0[246], M0[174], M0[143], M0[65], M0[48]};
layer0_N147 layer0_N147_inst (.M0(layer0_N147_wire), .M1(M1[295:294]));

wire [5:0] layer0_N148_wire = {M0[400], M0[327], M0[288], M0[215], M0[164], M0[92]};
layer0_N148 layer0_N148_inst (.M0(layer0_N148_wire), .M1(M1[297:296]));

wire [5:0] layer0_N149_wire = {M0[450], M0[409], M0[337], M0[334], M0[259], M0[25]};
layer0_N149 layer0_N149_inst (.M0(layer0_N149_wire), .M1(M1[299:298]));

wire [5:0] layer0_N150_wire = {M0[389], M0[322], M0[254], M0[248], M0[67], M0[38]};
layer0_N150 layer0_N150_inst (.M0(layer0_N150_wire), .M1(M1[301:300]));

wire [5:0] layer0_N151_wire = {M0[439], M0[407], M0[338], M0[309], M0[244], M0[53]};
layer0_N151 layer0_N151_inst (.M0(layer0_N151_wire), .M1(M1[303:302]));

wire [5:0] layer0_N152_wire = {M0[473], M0[451], M0[409], M0[347], M0[196], M0[65]};
layer0_N152 layer0_N152_inst (.M0(layer0_N152_wire), .M1(M1[305:304]));

wire [5:0] layer0_N153_wire = {M0[482], M0[440], M0[372], M0[316], M0[111], M0[74]};
layer0_N153 layer0_N153_inst (.M0(layer0_N153_wire), .M1(M1[307:306]));

wire [5:0] layer0_N154_wire = {M0[476], M0[355], M0[326], M0[172], M0[92], M0[84]};
layer0_N154 layer0_N154_inst (.M0(layer0_N154_wire), .M1(M1[309:308]));

wire [5:0] layer0_N155_wire = {M0[461], M0[359], M0[175], M0[157], M0[124], M0[26]};
layer0_N155 layer0_N155_inst (.M0(layer0_N155_wire), .M1(M1[311:310]));

wire [5:0] layer0_N156_wire = {M0[439], M0[247], M0[163], M0[161], M0[155], M0[138]};
layer0_N156 layer0_N156_inst (.M0(layer0_N156_wire), .M1(M1[313:312]));

wire [5:0] layer0_N157_wire = {M0[504], M0[110], M0[19], M0[16], M0[7], M0[5]};
layer0_N157 layer0_N157_inst (.M0(layer0_N157_wire), .M1(M1[315:314]));

wire [5:0] layer0_N158_wire = {M0[391], M0[339], M0[288], M0[230], M0[87], M0[49]};
layer0_N158 layer0_N158_inst (.M0(layer0_N158_wire), .M1(M1[317:316]));

wire [5:0] layer0_N159_wire = {M0[436], M0[427], M0[294], M0[246], M0[77], M0[27]};
layer0_N159 layer0_N159_inst (.M0(layer0_N159_wire), .M1(M1[319:318]));

wire [5:0] layer0_N160_wire = {M0[484], M0[442], M0[192], M0[129], M0[110], M0[109]};
layer0_N160 layer0_N160_inst (.M0(layer0_N160_wire), .M1(M1[321:320]));

wire [5:0] layer0_N161_wire = {M0[379], M0[369], M0[264], M0[244], M0[101], M0[94]};
layer0_N161 layer0_N161_inst (.M0(layer0_N161_wire), .M1(M1[323:322]));

wire [5:0] layer0_N162_wire = {M0[478], M0[440], M0[435], M0[180], M0[177], M0[62]};
layer0_N162 layer0_N162_inst (.M0(layer0_N162_wire), .M1(M1[325:324]));

wire [5:0] layer0_N163_wire = {M0[451], M0[384], M0[295], M0[130], M0[110], M0[78]};
layer0_N163 layer0_N163_inst (.M0(layer0_N163_wire), .M1(M1[327:326]));

wire [5:0] layer0_N164_wire = {M0[322], M0[307], M0[265], M0[249], M0[110], M0[26]};
layer0_N164 layer0_N164_inst (.M0(layer0_N164_wire), .M1(M1[329:328]));

wire [5:0] layer0_N165_wire = {M0[505], M0[495], M0[353], M0[278], M0[257], M0[186]};
layer0_N165 layer0_N165_inst (.M0(layer0_N165_wire), .M1(M1[331:330]));

wire [5:0] layer0_N166_wire = {M0[381], M0[182], M0[177], M0[131], M0[93], M0[65]};
layer0_N166 layer0_N166_inst (.M0(layer0_N166_wire), .M1(M1[333:332]));

wire [5:0] layer0_N167_wire = {M0[335], M0[208], M0[182], M0[142], M0[107], M0[59]};
layer0_N167 layer0_N167_inst (.M0(layer0_N167_wire), .M1(M1[335:334]));

wire [5:0] layer0_N168_wire = {M0[414], M0[291], M0[243], M0[196], M0[190], M0[96]};
layer0_N168 layer0_N168_inst (.M0(layer0_N168_wire), .M1(M1[337:336]));

wire [5:0] layer0_N169_wire = {M0[412], M0[340], M0[316], M0[264], M0[150], M0[25]};
layer0_N169 layer0_N169_inst (.M0(layer0_N169_wire), .M1(M1[339:338]));

wire [5:0] layer0_N170_wire = {M0[500], M0[456], M0[207], M0[101], M0[46], M0[24]};
layer0_N170 layer0_N170_inst (.M0(layer0_N170_wire), .M1(M1[341:340]));

wire [5:0] layer0_N171_wire = {M0[493], M0[374], M0[300], M0[294], M0[281], M0[86]};
layer0_N171 layer0_N171_inst (.M0(layer0_N171_wire), .M1(M1[343:342]));

wire [5:0] layer0_N172_wire = {M0[339], M0[298], M0[168], M0[89], M0[84], M0[48]};
layer0_N172 layer0_N172_inst (.M0(layer0_N172_wire), .M1(M1[345:344]));

wire [5:0] layer0_N173_wire = {M0[464], M0[463], M0[432], M0[255], M0[190], M0[73]};
layer0_N173 layer0_N173_inst (.M0(layer0_N173_wire), .M1(M1[347:346]));

wire [5:0] layer0_N174_wire = {M0[466], M0[359], M0[351], M0[325], M0[295], M0[211]};
layer0_N174 layer0_N174_inst (.M0(layer0_N174_wire), .M1(M1[349:348]));

wire [5:0] layer0_N175_wire = {M0[319], M0[233], M0[209], M0[156], M0[106], M0[23]};
layer0_N175 layer0_N175_inst (.M0(layer0_N175_wire), .M1(M1[351:350]));

wire [5:0] layer0_N176_wire = {M0[505], M0[446], M0[252], M0[241], M0[224], M0[8]};
layer0_N176 layer0_N176_inst (.M0(layer0_N176_wire), .M1(M1[353:352]));

wire [5:0] layer0_N177_wire = {M0[439], M0[436], M0[401], M0[380], M0[362], M0[116]};
layer0_N177 layer0_N177_inst (.M0(layer0_N177_wire), .M1(M1[355:354]));

wire [5:0] layer0_N178_wire = {M0[219], M0[143], M0[122], M0[54], M0[13], M0[4]};
layer0_N178 layer0_N178_inst (.M0(layer0_N178_wire), .M1(M1[357:356]));

wire [5:0] layer0_N179_wire = {M0[488], M0[380], M0[294], M0[241], M0[214], M0[21]};
layer0_N179 layer0_N179_inst (.M0(layer0_N179_wire), .M1(M1[359:358]));

wire [5:0] layer0_N180_wire = {M0[509], M0[472], M0[447], M0[313], M0[207], M0[32]};
layer0_N180 layer0_N180_inst (.M0(layer0_N180_wire), .M1(M1[361:360]));

wire [5:0] layer0_N181_wire = {M0[440], M0[212], M0[177], M0[167], M0[165], M0[163]};
layer0_N181 layer0_N181_inst (.M0(layer0_N181_wire), .M1(M1[363:362]));

wire [5:0] layer0_N182_wire = {M0[493], M0[349], M0[310], M0[288], M0[138], M0[8]};
layer0_N182 layer0_N182_inst (.M0(layer0_N182_wire), .M1(M1[365:364]));

wire [5:0] layer0_N183_wire = {M0[506], M0[474], M0[443], M0[408], M0[349], M0[308]};
layer0_N183 layer0_N183_inst (.M0(layer0_N183_wire), .M1(M1[367:366]));

wire [5:0] layer0_N184_wire = {M0[467], M0[433], M0[357], M0[268], M0[210], M0[205]};
layer0_N184 layer0_N184_inst (.M0(layer0_N184_wire), .M1(M1[369:368]));

wire [5:0] layer0_N185_wire = {M0[395], M0[328], M0[261], M0[210], M0[15], M0[2]};
layer0_N185 layer0_N185_inst (.M0(layer0_N185_wire), .M1(M1[371:370]));

wire [5:0] layer0_N186_wire = {M0[460], M0[454], M0[325], M0[304], M0[163], M0[101]};
layer0_N186 layer0_N186_inst (.M0(layer0_N186_wire), .M1(M1[373:372]));

wire [5:0] layer0_N187_wire = {M0[500], M0[449], M0[426], M0[377], M0[83], M0[76]};
layer0_N187 layer0_N187_inst (.M0(layer0_N187_wire), .M1(M1[375:374]));

wire [5:0] layer0_N188_wire = {M0[242], M0[201], M0[125], M0[27], M0[23], M0[1]};
layer0_N188 layer0_N188_inst (.M0(layer0_N188_wire), .M1(M1[377:376]));

wire [5:0] layer0_N189_wire = {M0[452], M0[288], M0[282], M0[190], M0[146], M0[124]};
layer0_N189 layer0_N189_inst (.M0(layer0_N189_wire), .M1(M1[379:378]));

wire [5:0] layer0_N190_wire = {M0[506], M0[485], M0[482], M0[435], M0[99], M0[26]};
layer0_N190 layer0_N190_inst (.M0(layer0_N190_wire), .M1(M1[381:380]));

wire [5:0] layer0_N191_wire = {M0[487], M0[474], M0[454], M0[428], M0[300], M0[13]};
layer0_N191 layer0_N191_inst (.M0(layer0_N191_wire), .M1(M1[383:382]));

wire [5:0] layer0_N192_wire = {M0[379], M0[342], M0[190], M0[189], M0[61], M0[1]};
layer0_N192 layer0_N192_inst (.M0(layer0_N192_wire), .M1(M1[385:384]));

wire [5:0] layer0_N193_wire = {M0[452], M0[403], M0[308], M0[279], M0[160], M0[77]};
layer0_N193 layer0_N193_inst (.M0(layer0_N193_wire), .M1(M1[387:386]));

wire [5:0] layer0_N194_wire = {M0[480], M0[471], M0[362], M0[329], M0[254], M0[177]};
layer0_N194 layer0_N194_inst (.M0(layer0_N194_wire), .M1(M1[389:388]));

wire [5:0] layer0_N195_wire = {M0[487], M0[158], M0[145], M0[54], M0[36], M0[29]};
layer0_N195 layer0_N195_inst (.M0(layer0_N195_wire), .M1(M1[391:390]));

wire [5:0] layer0_N196_wire = {M0[384], M0[214], M0[174], M0[120], M0[21], M0[4]};
layer0_N196 layer0_N196_inst (.M0(layer0_N196_wire), .M1(M1[393:392]));

wire [5:0] layer0_N197_wire = {M0[364], M0[362], M0[332], M0[308], M0[86], M0[58]};
layer0_N197 layer0_N197_inst (.M0(layer0_N197_wire), .M1(M1[395:394]));

wire [5:0] layer0_N198_wire = {M0[431], M0[397], M0[386], M0[269], M0[241], M0[186]};
layer0_N198 layer0_N198_inst (.M0(layer0_N198_wire), .M1(M1[397:396]));

wire [5:0] layer0_N199_wire = {M0[496], M0[449], M0[404], M0[351], M0[205], M0[60]};
layer0_N199 layer0_N199_inst (.M0(layer0_N199_wire), .M1(M1[399:398]));

wire [5:0] layer0_N200_wire = {M0[368], M0[323], M0[271], M0[262], M0[110], M0[74]};
layer0_N200 layer0_N200_inst (.M0(layer0_N200_wire), .M1(M1[401:400]));

wire [5:0] layer0_N201_wire = {M0[317], M0[306], M0[275], M0[63], M0[36], M0[24]};
layer0_N201 layer0_N201_inst (.M0(layer0_N201_wire), .M1(M1[403:402]));

wire [5:0] layer0_N202_wire = {M0[479], M0[451], M0[365], M0[226], M0[102], M0[18]};
layer0_N202 layer0_N202_inst (.M0(layer0_N202_wire), .M1(M1[405:404]));

wire [5:0] layer0_N203_wire = {M0[430], M0[393], M0[280], M0[196], M0[50], M0[7]};
layer0_N203 layer0_N203_inst (.M0(layer0_N203_wire), .M1(M1[407:406]));

wire [5:0] layer0_N204_wire = {M0[335], M0[222], M0[178], M0[164], M0[118], M0[67]};
layer0_N204 layer0_N204_inst (.M0(layer0_N204_wire), .M1(M1[409:408]));

wire [5:0] layer0_N205_wire = {M0[496], M0[475], M0[463], M0[223], M0[91], M0[69]};
layer0_N205 layer0_N205_inst (.M0(layer0_N205_wire), .M1(M1[411:410]));

wire [5:0] layer0_N206_wire = {M0[413], M0[412], M0[297], M0[268], M0[267], M0[67]};
layer0_N206 layer0_N206_inst (.M0(layer0_N206_wire), .M1(M1[413:412]));

wire [5:0] layer0_N207_wire = {M0[309], M0[285], M0[164], M0[140], M0[123], M0[103]};
layer0_N207 layer0_N207_inst (.M0(layer0_N207_wire), .M1(M1[415:414]));

wire [5:0] layer0_N208_wire = {M0[395], M0[316], M0[53], M0[26], M0[22], M0[18]};
layer0_N208 layer0_N208_inst (.M0(layer0_N208_wire), .M1(M1[417:416]));

wire [5:0] layer0_N209_wire = {M0[484], M0[385], M0[276], M0[230], M0[130], M0[100]};
layer0_N209 layer0_N209_inst (.M0(layer0_N209_wire), .M1(M1[419:418]));

wire [5:0] layer0_N210_wire = {M0[393], M0[337], M0[327], M0[321], M0[314], M0[294]};
layer0_N210 layer0_N210_inst (.M0(layer0_N210_wire), .M1(M1[421:420]));

wire [5:0] layer0_N211_wire = {M0[459], M0[394], M0[179], M0[150], M0[60], M0[12]};
layer0_N211 layer0_N211_inst (.M0(layer0_N211_wire), .M1(M1[423:422]));

wire [5:0] layer0_N212_wire = {M0[493], M0[488], M0[350], M0[265], M0[188], M0[181]};
layer0_N212 layer0_N212_inst (.M0(layer0_N212_wire), .M1(M1[425:424]));

wire [5:0] layer0_N213_wire = {M0[364], M0[353], M0[352], M0[199], M0[181], M0[92]};
layer0_N213 layer0_N213_inst (.M0(layer0_N213_wire), .M1(M1[427:426]));

wire [5:0] layer0_N214_wire = {M0[488], M0[289], M0[285], M0[258], M0[152], M0[94]};
layer0_N214 layer0_N214_inst (.M0(layer0_N214_wire), .M1(M1[429:428]));

wire [5:0] layer0_N215_wire = {M0[484], M0[373], M0[355], M0[241], M0[166], M0[0]};
layer0_N215 layer0_N215_inst (.M0(layer0_N215_wire), .M1(M1[431:430]));

wire [5:0] layer0_N216_wire = {M0[313], M0[210], M0[185], M0[64], M0[48], M0[16]};
layer0_N216 layer0_N216_inst (.M0(layer0_N216_wire), .M1(M1[433:432]));

wire [5:0] layer0_N217_wire = {M0[331], M0[104], M0[78], M0[63], M0[43], M0[31]};
layer0_N217 layer0_N217_inst (.M0(layer0_N217_wire), .M1(M1[435:434]));

wire [5:0] layer0_N218_wire = {M0[443], M0[428], M0[418], M0[412], M0[209], M0[44]};
layer0_N218 layer0_N218_inst (.M0(layer0_N218_wire), .M1(M1[437:436]));

wire [5:0] layer0_N219_wire = {M0[491], M0[283], M0[182], M0[176], M0[142], M0[7]};
layer0_N219 layer0_N219_inst (.M0(layer0_N219_wire), .M1(M1[439:438]));

wire [5:0] layer0_N220_wire = {M0[459], M0[380], M0[278], M0[184], M0[77], M0[67]};
layer0_N220 layer0_N220_inst (.M0(layer0_N220_wire), .M1(M1[441:440]));

wire [5:0] layer0_N221_wire = {M0[475], M0[347], M0[338], M0[309], M0[144], M0[40]};
layer0_N221 layer0_N221_inst (.M0(layer0_N221_wire), .M1(M1[443:442]));

wire [5:0] layer0_N222_wire = {M0[506], M0[226], M0[176], M0[120], M0[65], M0[52]};
layer0_N222 layer0_N222_inst (.M0(layer0_N222_wire), .M1(M1[445:444]));

wire [5:0] layer0_N223_wire = {M0[398], M0[260], M0[199], M0[179], M0[94], M0[41]};
layer0_N223 layer0_N223_inst (.M0(layer0_N223_wire), .M1(M1[447:446]));

wire [5:0] layer0_N224_wire = {M0[418], M0[351], M0[218], M0[123], M0[49], M0[2]};
layer0_N224 layer0_N224_inst (.M0(layer0_N224_wire), .M1(M1[449:448]));

wire [5:0] layer0_N225_wire = {M0[371], M0[313], M0[281], M0[221], M0[142], M0[47]};
layer0_N225 layer0_N225_inst (.M0(layer0_N225_wire), .M1(M1[451:450]));

wire [5:0] layer0_N226_wire = {M0[401], M0[369], M0[267], M0[164], M0[53], M0[23]};
layer0_N226 layer0_N226_inst (.M0(layer0_N226_wire), .M1(M1[453:452]));

wire [5:0] layer0_N227_wire = {M0[486], M0[410], M0[397], M0[357], M0[190], M0[48]};
layer0_N227 layer0_N227_inst (.M0(layer0_N227_wire), .M1(M1[455:454]));

wire [5:0] layer0_N228_wire = {M0[351], M0[342], M0[304], M0[270], M0[11], M0[4]};
layer0_N228 layer0_N228_inst (.M0(layer0_N228_wire), .M1(M1[457:456]));

wire [5:0] layer0_N229_wire = {M0[493], M0[166], M0[133], M0[131], M0[120], M0[75]};
layer0_N229 layer0_N229_inst (.M0(layer0_N229_wire), .M1(M1[459:458]));

wire [5:0] layer0_N230_wire = {M0[391], M0[356], M0[237], M0[48], M0[27], M0[6]};
layer0_N230 layer0_N230_inst (.M0(layer0_N230_wire), .M1(M1[461:460]));

wire [5:0] layer0_N231_wire = {M0[204], M0[199], M0[189], M0[155], M0[149], M0[20]};
layer0_N231 layer0_N231_inst (.M0(layer0_N231_wire), .M1(M1[463:462]));

wire [5:0] layer0_N232_wire = {M0[450], M0[346], M0[314], M0[202], M0[189], M0[25]};
layer0_N232 layer0_N232_inst (.M0(layer0_N232_wire), .M1(M1[465:464]));

wire [5:0] layer0_N233_wire = {M0[503], M0[502], M0[154], M0[25], M0[23], M0[21]};
layer0_N233 layer0_N233_inst (.M0(layer0_N233_wire), .M1(M1[467:466]));

wire [5:0] layer0_N234_wire = {M0[492], M0[454], M0[341], M0[312], M0[197], M0[86]};
layer0_N234 layer0_N234_inst (.M0(layer0_N234_wire), .M1(M1[469:468]));

wire [5:0] layer0_N235_wire = {M0[435], M0[313], M0[305], M0[290], M0[186], M0[56]};
layer0_N235 layer0_N235_inst (.M0(layer0_N235_wire), .M1(M1[471:470]));

wire [5:0] layer0_N236_wire = {M0[509], M0[491], M0[429], M0[375], M0[292], M0[120]};
layer0_N236 layer0_N236_inst (.M0(layer0_N236_wire), .M1(M1[473:472]));

wire [5:0] layer0_N237_wire = {M0[426], M0[296], M0[248], M0[63], M0[61], M0[33]};
layer0_N237 layer0_N237_inst (.M0(layer0_N237_wire), .M1(M1[475:474]));

wire [5:0] layer0_N238_wire = {M0[415], M0[336], M0[310], M0[213], M0[165], M0[160]};
layer0_N238 layer0_N238_inst (.M0(layer0_N238_wire), .M1(M1[477:476]));

wire [5:0] layer0_N239_wire = {M0[471], M0[265], M0[253], M0[210], M0[199], M0[102]};
layer0_N239 layer0_N239_inst (.M0(layer0_N239_wire), .M1(M1[479:478]));

wire [5:0] layer0_N240_wire = {M0[405], M0[341], M0[307], M0[153], M0[129], M0[31]};
layer0_N240 layer0_N240_inst (.M0(layer0_N240_wire), .M1(M1[481:480]));

wire [5:0] layer0_N241_wire = {M0[398], M0[317], M0[152], M0[113], M0[102], M0[70]};
layer0_N241 layer0_N241_inst (.M0(layer0_N241_wire), .M1(M1[483:482]));

wire [5:0] layer0_N242_wire = {M0[355], M0[306], M0[265], M0[229], M0[219], M0[24]};
layer0_N242 layer0_N242_inst (.M0(layer0_N242_wire), .M1(M1[485:484]));

wire [5:0] layer0_N243_wire = {M0[434], M0[250], M0[221], M0[152], M0[79], M0[1]};
layer0_N243 layer0_N243_inst (.M0(layer0_N243_wire), .M1(M1[487:486]));

wire [5:0] layer0_N244_wire = {M0[499], M0[489], M0[383], M0[377], M0[355], M0[93]};
layer0_N244 layer0_N244_inst (.M0(layer0_N244_wire), .M1(M1[489:488]));

wire [5:0] layer0_N245_wire = {M0[503], M0[406], M0[362], M0[317], M0[220], M0[121]};
layer0_N245 layer0_N245_inst (.M0(layer0_N245_wire), .M1(M1[491:490]));

wire [5:0] layer0_N246_wire = {M0[422], M0[376], M0[354], M0[292], M0[73], M0[66]};
layer0_N246 layer0_N246_inst (.M0(layer0_N246_wire), .M1(M1[493:492]));

wire [5:0] layer0_N247_wire = {M0[494], M0[424], M0[87], M0[43], M0[39], M0[7]};
layer0_N247 layer0_N247_inst (.M0(layer0_N247_wire), .M1(M1[495:494]));

wire [5:0] layer0_N248_wire = {M0[332], M0[326], M0[268], M0[242], M0[156], M0[21]};
layer0_N248 layer0_N248_inst (.M0(layer0_N248_wire), .M1(M1[497:496]));

wire [5:0] layer0_N249_wire = {M0[498], M0[434], M0[383], M0[374], M0[264], M0[51]};
layer0_N249 layer0_N249_inst (.M0(layer0_N249_wire), .M1(M1[499:498]));

wire [5:0] layer0_N250_wire = {M0[357], M0[217], M0[162], M0[104], M0[51], M0[12]};
layer0_N250 layer0_N250_inst (.M0(layer0_N250_wire), .M1(M1[501:500]));

wire [5:0] layer0_N251_wire = {M0[403], M0[369], M0[311], M0[121], M0[94], M0[68]};
layer0_N251 layer0_N251_inst (.M0(layer0_N251_wire), .M1(M1[503:502]));

wire [5:0] layer0_N252_wire = {M0[389], M0[168], M0[155], M0[134], M0[116], M0[41]};
layer0_N252 layer0_N252_inst (.M0(layer0_N252_wire), .M1(M1[505:504]));

wire [5:0] layer0_N253_wire = {M0[485], M0[468], M0[464], M0[293], M0[140], M0[58]};
layer0_N253 layer0_N253_inst (.M0(layer0_N253_wire), .M1(M1[507:506]));

wire [5:0] layer0_N254_wire = {M0[389], M0[210], M0[195], M0[60], M0[11], M0[2]};
layer0_N254 layer0_N254_inst (.M0(layer0_N254_wire), .M1(M1[509:508]));

wire [5:0] layer0_N255_wire = {M0[464], M0[364], M0[345], M0[272], M0[165], M0[128]};
layer0_N255 layer0_N255_inst (.M0(layer0_N255_wire), .M1(M1[511:510]));

endmodule