module layer1 (input [1185:0] M0, output [199:0] M1);

wire [5:0] layer1_N0_wire = {M0[385], M0[384], M0[111], M0[110], M0[93], M0[92]};
layer1_N0 layer1_N0_inst (.M0(layer1_N0_wire), .M1(M1[1:0]));

wire [5:0] layer1_N1_wire = {M0[439], M0[438], M0[429], M0[428], M0[299], M0[298]};
layer1_N1 layer1_N1_inst (.M0(layer1_N1_wire), .M1(M1[3:2]));

wire [5:0] layer1_N2_wire = {M0[775], M0[774], M0[535], M0[534], M0[205], M0[204]};
layer1_N2 layer1_N2_inst (.M0(layer1_N2_wire), .M1(M1[5:4]));

wire [5:0] layer1_N3_wire = {M0[703], M0[702], M0[161], M0[160], M0[157], M0[156]};
layer1_N3 layer1_N3_inst (.M0(layer1_N3_wire), .M1(M1[7:6]));

wire [5:0] layer1_N4_wire = {M0[517], M0[516], M0[411], M0[410], M0[65], M0[64]};
layer1_N4 layer1_N4_inst (.M0(layer1_N4_wire), .M1(M1[9:8]));

wire [5:0] layer1_N5_wire = {M0[1039], M0[1038], M0[705], M0[704], M0[435], M0[434]};
layer1_N5 layer1_N5_inst (.M0(layer1_N5_wire), .M1(M1[11:10]));

wire [5:0] layer1_N6_wire = {M0[851], M0[850], M0[717], M0[716], M0[693], M0[692]};
layer1_N6 layer1_N6_inst (.M0(layer1_N6_wire), .M1(M1[13:12]));

wire [5:0] layer1_N7_wire = {M0[871], M0[870], M0[511], M0[510], M0[397], M0[396]};
layer1_N7 layer1_N7_inst (.M0(layer1_N7_wire), .M1(M1[15:14]));

wire [5:0] layer1_N8_wire = {M0[919], M0[918], M0[383], M0[382], M0[99], M0[98]};
layer1_N8 layer1_N8_inst (.M0(layer1_N8_wire), .M1(M1[17:16]));

wire [5:0] layer1_N9_wire = {M0[1091], M0[1090], M0[753], M0[752], M0[579], M0[578]};
layer1_N9 layer1_N9_inst (.M0(layer1_N9_wire), .M1(M1[19:18]));

wire [5:0] layer1_N10_wire = {M0[601], M0[600], M0[549], M0[548], M0[441], M0[440]};
layer1_N10 layer1_N10_inst (.M0(layer1_N10_wire), .M1(M1[21:20]));

wire [5:0] layer1_N11_wire = {M0[837], M0[836], M0[655], M0[654], M0[265], M0[264]};
layer1_N11 layer1_N11_inst (.M0(layer1_N11_wire), .M1(M1[23:22]));

wire [5:0] layer1_N12_wire = {M0[1119], M0[1118], M0[325], M0[324], M0[29], M0[28]};
layer1_N12 layer1_N12_inst (.M0(layer1_N12_wire), .M1(M1[25:24]));

wire [5:0] layer1_N13_wire = {M0[835], M0[834], M0[437], M0[436], M0[203], M0[202]};
layer1_N13 layer1_N13_inst (.M0(layer1_N13_wire), .M1(M1[27:26]));

wire [5:0] layer1_N14_wire = {M0[693], M0[692], M0[215], M0[214], M0[19], M0[18]};
layer1_N14 layer1_N14_inst (.M0(layer1_N14_wire), .M1(M1[29:28]));

wire [5:0] layer1_N15_wire = {M0[871], M0[870], M0[815], M0[814], M0[557], M0[556]};
layer1_N15 layer1_N15_inst (.M0(layer1_N15_wire), .M1(M1[31:30]));

wire [5:0] layer1_N16_wire = {M0[965], M0[964], M0[591], M0[590], M0[251], M0[250]};
layer1_N16 layer1_N16_inst (.M0(layer1_N16_wire), .M1(M1[33:32]));

wire [5:0] layer1_N17_wire = {M0[883], M0[882], M0[627], M0[626], M0[327], M0[326]};
layer1_N17 layer1_N17_inst (.M0(layer1_N17_wire), .M1(M1[35:34]));

wire [5:0] layer1_N18_wire = {M0[795], M0[794], M0[761], M0[760], M0[603], M0[602]};
layer1_N18 layer1_N18_inst (.M0(layer1_N18_wire), .M1(M1[37:36]));

wire [5:0] layer1_N19_wire = {M0[771], M0[770], M0[525], M0[524], M0[303], M0[302]};
layer1_N19 layer1_N19_inst (.M0(layer1_N19_wire), .M1(M1[39:38]));

wire [5:0] layer1_N20_wire = {M0[983], M0[982], M0[799], M0[798], M0[425], M0[424]};
layer1_N20 layer1_N20_inst (.M0(layer1_N20_wire), .M1(M1[41:40]));

wire [5:0] layer1_N21_wire = {M0[1155], M0[1154], M0[359], M0[358], M0[259], M0[258]};
layer1_N21 layer1_N21_inst (.M0(layer1_N21_wire), .M1(M1[43:42]));

wire [5:0] layer1_N22_wire = {M0[1125], M0[1124], M0[807], M0[806], M0[333], M0[332]};
layer1_N22 layer1_N22_inst (.M0(layer1_N22_wire), .M1(M1[45:44]));

wire [5:0] layer1_N23_wire = {M0[885], M0[884], M0[193], M0[192], M0[81], M0[80]};
layer1_N23 layer1_N23_inst (.M0(layer1_N23_wire), .M1(M1[47:46]));

wire [5:0] layer1_N24_wire = {M0[1153], M0[1152], M0[395], M0[394], M0[391], M0[390]};
layer1_N24 layer1_N24_inst (.M0(layer1_N24_wire), .M1(M1[49:48]));

wire [5:0] layer1_N25_wire = {M0[1137], M0[1136], M0[261], M0[260], M0[149], M0[148]};
layer1_N25 layer1_N25_inst (.M0(layer1_N25_wire), .M1(M1[51:50]));

wire [5:0] layer1_N26_wire = {M0[879], M0[878], M0[837], M0[836], M0[729], M0[728]};
layer1_N26 layer1_N26_inst (.M0(layer1_N26_wire), .M1(M1[53:52]));

wire [5:0] layer1_N27_wire = {M0[1067], M0[1066], M0[715], M0[714], M0[317], M0[316]};
layer1_N27 layer1_N27_inst (.M0(layer1_N27_wire), .M1(M1[55:54]));

wire [5:0] layer1_N28_wire = {M0[1019], M0[1018], M0[725], M0[724], M0[557], M0[556]};
layer1_N28 layer1_N28_inst (.M0(layer1_N28_wire), .M1(M1[57:56]));

wire [5:0] layer1_N29_wire = {M0[463], M0[462], M0[163], M0[162], M0[15], M0[14]};
layer1_N29 layer1_N29_inst (.M0(layer1_N29_wire), .M1(M1[59:58]));

wire [5:0] layer1_N30_wire = {M0[563], M0[562], M0[423], M0[422], M0[21], M0[20]};
layer1_N30 layer1_N30_inst (.M0(layer1_N30_wire), .M1(M1[61:60]));

wire [5:0] layer1_N31_wire = {M0[895], M0[894], M0[765], M0[764], M0[161], M0[160]};
layer1_N31 layer1_N31_inst (.M0(layer1_N31_wire), .M1(M1[63:62]));

wire [5:0] layer1_N32_wire = {M0[921], M0[920], M0[761], M0[760], M0[35], M0[34]};
layer1_N32 layer1_N32_inst (.M0(layer1_N32_wire), .M1(M1[65:64]));

wire [5:0] layer1_N33_wire = {M0[1177], M0[1176], M0[257], M0[256], M0[59], M0[58]};
layer1_N33 layer1_N33_inst (.M0(layer1_N33_wire), .M1(M1[67:66]));

wire [5:0] layer1_N34_wire = {M0[831], M0[830], M0[721], M0[720], M0[445], M0[444]};
layer1_N34 layer1_N34_inst (.M0(layer1_N34_wire), .M1(M1[69:68]));

wire [5:0] layer1_N35_wire = {M0[1147], M0[1146], M0[1027], M0[1026], M0[445], M0[444]};
layer1_N35 layer1_N35_inst (.M0(layer1_N35_wire), .M1(M1[71:70]));

wire [5:0] layer1_N36_wire = {M0[1035], M0[1034], M0[965], M0[964], M0[473], M0[472]};
layer1_N36 layer1_N36_inst (.M0(layer1_N36_wire), .M1(M1[73:72]));

wire [5:0] layer1_N37_wire = {M0[1007], M0[1006], M0[627], M0[626], M0[129], M0[128]};
layer1_N37 layer1_N37_inst (.M0(layer1_N37_wire), .M1(M1[75:74]));

wire [5:0] layer1_N38_wire = {M0[1139], M0[1138], M0[261], M0[260], M0[165], M0[164]};
layer1_N38 layer1_N38_inst (.M0(layer1_N38_wire), .M1(M1[77:76]));

wire [5:0] layer1_N39_wire = {M0[793], M0[792], M0[641], M0[640], M0[21], M0[20]};
layer1_N39 layer1_N39_inst (.M0(layer1_N39_wire), .M1(M1[79:78]));

wire [5:0] layer1_N40_wire = {M0[1041], M0[1040], M0[631], M0[630], M0[73], M0[72]};
layer1_N40 layer1_N40_inst (.M0(layer1_N40_wire), .M1(M1[81:80]));

wire [5:0] layer1_N41_wire = {M0[1173], M0[1172], M0[1017], M0[1016], M0[727], M0[726]};
layer1_N41 layer1_N41_inst (.M0(layer1_N41_wire), .M1(M1[83:82]));

wire [5:0] layer1_N42_wire = {M0[355], M0[354], M0[133], M0[132], M0[79], M0[78]};
layer1_N42 layer1_N42_inst (.M0(layer1_N42_wire), .M1(M1[85:84]));

wire [5:0] layer1_N43_wire = {M0[1181], M0[1180], M0[1065], M0[1064], M0[593], M0[592]};
layer1_N43 layer1_N43_inst (.M0(layer1_N43_wire), .M1(M1[87:86]));

wire [5:0] layer1_N44_wire = {M0[873], M0[872], M0[645], M0[644], M0[211], M0[210]};
layer1_N44 layer1_N44_inst (.M0(layer1_N44_wire), .M1(M1[89:88]));

wire [5:0] layer1_N45_wire = {M0[1179], M0[1178], M0[647], M0[646], M0[327], M0[326]};
layer1_N45 layer1_N45_inst (.M0(layer1_N45_wire), .M1(M1[91:90]));

wire [5:0] layer1_N46_wire = {M0[1089], M0[1088], M0[287], M0[286], M0[129], M0[128]};
layer1_N46 layer1_N46_inst (.M0(layer1_N46_wire), .M1(M1[93:92]));

wire [5:0] layer1_N47_wire = {M0[863], M0[862], M0[805], M0[804], M0[167], M0[166]};
layer1_N47 layer1_N47_inst (.M0(layer1_N47_wire), .M1(M1[95:94]));

wire [5:0] layer1_N48_wire = {M0[1039], M0[1038], M0[859], M0[858], M0[337], M0[336]};
layer1_N48 layer1_N48_inst (.M0(layer1_N48_wire), .M1(M1[97:96]));

wire [5:0] layer1_N49_wire = {M0[491], M0[490], M0[221], M0[220], M0[13], M0[12]};
layer1_N49 layer1_N49_inst (.M0(layer1_N49_wire), .M1(M1[99:98]));

wire [5:0] layer1_N50_wire = {M0[1185], M0[1184], M0[173], M0[172], M0[111], M0[110]};
layer1_N50 layer1_N50_inst (.M0(layer1_N50_wire), .M1(M1[101:100]));

wire [5:0] layer1_N51_wire = {M0[769], M0[768], M0[425], M0[424], M0[59], M0[58]};
layer1_N51 layer1_N51_inst (.M0(layer1_N51_wire), .M1(M1[103:102]));

wire [5:0] layer1_N52_wire = {M0[1067], M0[1066], M0[1057], M0[1056], M0[771], M0[770]};
layer1_N52 layer1_N52_inst (.M0(layer1_N52_wire), .M1(M1[105:104]));

wire [5:0] layer1_N53_wire = {M0[1067], M0[1066], M0[927], M0[926], M0[497], M0[496]};
layer1_N53 layer1_N53_inst (.M0(layer1_N53_wire), .M1(M1[107:106]));

wire [5:0] layer1_N54_wire = {M0[1121], M0[1120], M0[763], M0[762], M0[405], M0[404]};
layer1_N54 layer1_N54_inst (.M0(layer1_N54_wire), .M1(M1[109:108]));

wire [5:0] layer1_N55_wire = {M0[1115], M0[1114], M0[629], M0[628], M0[199], M0[198]};
layer1_N55 layer1_N55_inst (.M0(layer1_N55_wire), .M1(M1[111:110]));

wire [5:0] layer1_N56_wire = {M0[703], M0[702], M0[517], M0[516], M0[31], M0[30]};
layer1_N56 layer1_N56_inst (.M0(layer1_N56_wire), .M1(M1[113:112]));

wire [5:0] layer1_N57_wire = {M0[1119], M0[1118], M0[691], M0[690], M0[221], M0[220]};
layer1_N57 layer1_N57_inst (.M0(layer1_N57_wire), .M1(M1[115:114]));

wire [5:0] layer1_N58_wire = {M0[1123], M0[1122], M0[1119], M0[1118], M0[905], M0[904]};
layer1_N58 layer1_N58_inst (.M0(layer1_N58_wire), .M1(M1[117:116]));

wire [5:0] layer1_N59_wire = {M0[781], M0[780], M0[461], M0[460], M0[433], M0[432]};
layer1_N59 layer1_N59_inst (.M0(layer1_N59_wire), .M1(M1[119:118]));

wire [5:0] layer1_N60_wire = {M0[1181], M0[1180], M0[1033], M0[1032], M0[491], M0[490]};
layer1_N60 layer1_N60_inst (.M0(layer1_N60_wire), .M1(M1[121:120]));

wire [5:0] layer1_N61_wire = {M0[879], M0[878], M0[229], M0[228], M0[183], M0[182]};
layer1_N61 layer1_N61_inst (.M0(layer1_N61_wire), .M1(M1[123:122]));

wire [5:0] layer1_N62_wire = {M0[1011], M0[1010], M0[699], M0[698], M0[61], M0[60]};
layer1_N62 layer1_N62_inst (.M0(layer1_N62_wire), .M1(M1[125:124]));

wire [5:0] layer1_N63_wire = {M0[903], M0[902], M0[585], M0[584], M0[135], M0[134]};
layer1_N63 layer1_N63_inst (.M0(layer1_N63_wire), .M1(M1[127:126]));

wire [5:0] layer1_N64_wire = {M0[775], M0[774], M0[419], M0[418], M0[121], M0[120]};
layer1_N64 layer1_N64_inst (.M0(layer1_N64_wire), .M1(M1[129:128]));

wire [5:0] layer1_N65_wire = {M0[1145], M0[1144], M0[917], M0[916], M0[543], M0[542]};
layer1_N65 layer1_N65_inst (.M0(layer1_N65_wire), .M1(M1[131:130]));

wire [5:0] layer1_N66_wire = {M0[871], M0[870], M0[139], M0[138], M0[39], M0[38]};
layer1_N66 layer1_N66_inst (.M0(layer1_N66_wire), .M1(M1[133:132]));

wire [5:0] layer1_N67_wire = {M0[1159], M0[1158], M0[1019], M0[1018], M0[153], M0[152]};
layer1_N67 layer1_N67_inst (.M0(layer1_N67_wire), .M1(M1[135:134]));

wire [5:0] layer1_N68_wire = {M0[1045], M0[1044], M0[979], M0[978], M0[37], M0[36]};
layer1_N68 layer1_N68_inst (.M0(layer1_N68_wire), .M1(M1[137:136]));

wire [5:0] layer1_N69_wire = {M0[1015], M0[1014], M0[963], M0[962], M0[397], M0[396]};
layer1_N69 layer1_N69_inst (.M0(layer1_N69_wire), .M1(M1[139:138]));

wire [5:0] layer1_N70_wire = {M0[443], M0[442], M0[343], M0[342], M0[53], M0[52]};
layer1_N70 layer1_N70_inst (.M0(layer1_N70_wire), .M1(M1[141:140]));

wire [5:0] layer1_N71_wire = {M0[1149], M0[1148], M0[555], M0[554], M0[399], M0[398]};
layer1_N71 layer1_N71_inst (.M0(layer1_N71_wire), .M1(M1[143:142]));

wire [5:0] layer1_N72_wire = {M0[1123], M0[1122], M0[1033], M0[1032], M0[961], M0[960]};
layer1_N72 layer1_N72_inst (.M0(layer1_N72_wire), .M1(M1[145:144]));

wire [5:0] layer1_N73_wire = {M0[1101], M0[1100], M0[757], M0[756], M0[105], M0[104]};
layer1_N73 layer1_N73_inst (.M0(layer1_N73_wire), .M1(M1[147:146]));

wire [5:0] layer1_N74_wire = {M0[783], M0[782], M0[629], M0[628], M0[321], M0[320]};
layer1_N74 layer1_N74_inst (.M0(layer1_N74_wire), .M1(M1[149:148]));

wire [5:0] layer1_N75_wire = {M0[1105], M0[1104], M0[109], M0[108], M0[69], M0[68]};
layer1_N75 layer1_N75_inst (.M0(layer1_N75_wire), .M1(M1[151:150]));

wire [5:0] layer1_N76_wire = {M0[951], M0[950], M0[897], M0[896], M0[609], M0[608]};
layer1_N76 layer1_N76_inst (.M0(layer1_N76_wire), .M1(M1[153:152]));

wire [5:0] layer1_N77_wire = {M0[1161], M0[1160], M0[183], M0[182], M0[73], M0[72]};
layer1_N77 layer1_N77_inst (.M0(layer1_N77_wire), .M1(M1[155:154]));

wire [5:0] layer1_N78_wire = {M0[1087], M0[1086], M0[985], M0[984], M0[479], M0[478]};
layer1_N78 layer1_N78_inst (.M0(layer1_N78_wire), .M1(M1[157:156]));

wire [5:0] layer1_N79_wire = {M0[753], M0[752], M0[553], M0[552], M0[55], M0[54]};
layer1_N79 layer1_N79_inst (.M0(layer1_N79_wire), .M1(M1[159:158]));

wire [5:0] layer1_N80_wire = {M0[775], M0[774], M0[705], M0[704], M0[265], M0[264]};
layer1_N80 layer1_N80_inst (.M0(layer1_N80_wire), .M1(M1[161:160]));

wire [5:0] layer1_N81_wire = {M0[887], M0[886], M0[867], M0[866], M0[809], M0[808]};
layer1_N81 layer1_N81_inst (.M0(layer1_N81_wire), .M1(M1[163:162]));

wire [5:0] layer1_N82_wire = {M0[1139], M0[1138], M0[1099], M0[1098], M0[845], M0[844]};
layer1_N82 layer1_N82_inst (.M0(layer1_N82_wire), .M1(M1[165:164]));

wire [5:0] layer1_N83_wire = {M0[529], M0[528], M0[375], M0[374], M0[367], M0[366]};
layer1_N83 layer1_N83_inst (.M0(layer1_N83_wire), .M1(M1[167:166]));

wire [5:0] layer1_N84_wire = {M0[791], M0[790], M0[767], M0[766], M0[469], M0[468]};
layer1_N84 layer1_N84_inst (.M0(layer1_N84_wire), .M1(M1[169:168]));

wire [5:0] layer1_N85_wire = {M0[1037], M0[1036], M0[623], M0[622], M0[415], M0[414]};
layer1_N85 layer1_N85_inst (.M0(layer1_N85_wire), .M1(M1[171:170]));

wire [5:0] layer1_N86_wire = {M0[1077], M0[1076], M0[309], M0[308], M0[305], M0[304]};
layer1_N86 layer1_N86_inst (.M0(layer1_N86_wire), .M1(M1[173:172]));

wire [5:0] layer1_N87_wire = {M0[877], M0[876], M0[479], M0[478], M0[99], M0[98]};
layer1_N87 layer1_N87_inst (.M0(layer1_N87_wire), .M1(M1[175:174]));

wire [5:0] layer1_N88_wire = {M0[749], M0[748], M0[575], M0[574], M0[269], M0[268]};
layer1_N88 layer1_N88_inst (.M0(layer1_N88_wire), .M1(M1[177:176]));

wire [5:0] layer1_N89_wire = {M0[721], M0[720], M0[713], M0[712], M0[573], M0[572]};
layer1_N89 layer1_N89_inst (.M0(layer1_N89_wire), .M1(M1[179:178]));

wire [5:0] layer1_N90_wire = {M0[951], M0[950], M0[917], M0[916], M0[809], M0[808]};
layer1_N90 layer1_N90_inst (.M0(layer1_N90_wire), .M1(M1[181:180]));

wire [5:0] layer1_N91_wire = {M0[953], M0[952], M0[453], M0[452], M0[11], M0[10]};
layer1_N91 layer1_N91_inst (.M0(layer1_N91_wire), .M1(M1[183:182]));

wire [5:0] layer1_N92_wire = {M0[1081], M0[1080], M0[849], M0[848], M0[669], M0[668]};
layer1_N92 layer1_N92_inst (.M0(layer1_N92_wire), .M1(M1[185:184]));

wire [5:0] layer1_N93_wire = {M0[977], M0[976], M0[251], M0[250], M0[235], M0[234]};
layer1_N93 layer1_N93_inst (.M0(layer1_N93_wire), .M1(M1[187:186]));

wire [5:0] layer1_N94_wire = {M0[1015], M0[1014], M0[711], M0[710], M0[475], M0[474]};
layer1_N94 layer1_N94_inst (.M0(layer1_N94_wire), .M1(M1[189:188]));

wire [5:0] layer1_N95_wire = {M0[1175], M0[1174], M0[935], M0[934], M0[429], M0[428]};
layer1_N95 layer1_N95_inst (.M0(layer1_N95_wire), .M1(M1[191:190]));

wire [5:0] layer1_N96_wire = {M0[599], M0[598], M0[473], M0[472], M0[225], M0[224]};
layer1_N96 layer1_N96_inst (.M0(layer1_N96_wire), .M1(M1[193:192]));

wire [5:0] layer1_N97_wire = {M0[1003], M0[1002], M0[203], M0[202], M0[5], M0[4]};
layer1_N97 layer1_N97_inst (.M0(layer1_N97_wire), .M1(M1[195:194]));

wire [5:0] layer1_N98_wire = {M0[669], M0[668], M0[449], M0[448], M0[391], M0[390]};
layer1_N98 layer1_N98_inst (.M0(layer1_N98_wire), .M1(M1[197:196]));

wire [5:0] layer1_N99_wire = {M0[975], M0[974], M0[93], M0[92], M0[51], M0[50]};
layer1_N99 layer1_N99_inst (.M0(layer1_N99_wire), .M1(M1[199:198]));

endmodule