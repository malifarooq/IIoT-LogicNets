module layer0 (input [511:0] M0, output [1185:0] M1);

wire [2:0] layer0_N0_wire = {M0[474], M0[353], M0[262]};
layer0_N0 layer0_N0_inst (.M0(layer0_N0_wire), .M1(M1[1:0]));

wire [2:0] layer0_N1_wire = {M0[436], M0[398], M0[270]};
layer0_N1 layer0_N1_inst (.M0(layer0_N1_wire), .M1(M1[3:2]));

wire [2:0] layer0_N2_wire = {M0[467], M0[143], M0[95]};
layer0_N2 layer0_N2_inst (.M0(layer0_N2_wire), .M1(M1[5:4]));

wire [2:0] layer0_N3_wire = {M0[500], M0[315], M0[220]};
layer0_N3 layer0_N3_inst (.M0(layer0_N3_wire), .M1(M1[7:6]));

wire [2:0] layer0_N4_wire = {M0[299], M0[20], M0[4]};
layer0_N4 layer0_N4_inst (.M0(layer0_N4_wire), .M1(M1[9:8]));

wire [2:0] layer0_N5_wire = {M0[388], M0[254], M0[48]};
layer0_N5 layer0_N5_inst (.M0(layer0_N5_wire), .M1(M1[11:10]));

wire [2:0] layer0_N6_wire = {M0[497], M0[494], M0[249]};
layer0_N6 layer0_N6_inst (.M0(layer0_N6_wire), .M1(M1[13:12]));

wire [2:0] layer0_N7_wire = {M0[356], M0[164], M0[142]};
layer0_N7 layer0_N7_inst (.M0(layer0_N7_wire), .M1(M1[15:14]));

wire [2:0] layer0_N8_wire = {M0[457], M0[382], M0[225]};
layer0_N8 layer0_N8_inst (.M0(layer0_N8_wire), .M1(M1[17:16]));

wire [2:0] layer0_N9_wire = {M0[472], M0[375], M0[14]};
layer0_N9 layer0_N9_inst (.M0(layer0_N9_wire), .M1(M1[19:18]));

wire [2:0] layer0_N10_wire = {M0[486], M0[410], M0[359]};
layer0_N10 layer0_N10_inst (.M0(layer0_N10_wire), .M1(M1[21:20]));

wire [2:0] layer0_N11_wire = {M0[372], M0[262], M0[151]};
layer0_N11 layer0_N11_inst (.M0(layer0_N11_wire), .M1(M1[23:22]));

wire [2:0] layer0_N12_wire = {M0[474], M0[284], M0[89]};
layer0_N12 layer0_N12_inst (.M0(layer0_N12_wire), .M1(M1[25:24]));

wire [2:0] layer0_N13_wire = {M0[427], M0[322], M0[136]};
layer0_N13 layer0_N13_inst (.M0(layer0_N13_wire), .M1(M1[27:26]));

wire [2:0] layer0_N14_wire = {M0[348], M0[154], M0[152]};
layer0_N14 layer0_N14_inst (.M0(layer0_N14_wire), .M1(M1[29:28]));

wire [2:0] layer0_N15_wire = {M0[409], M0[395], M0[152]};
layer0_N15 layer0_N15_inst (.M0(layer0_N15_wire), .M1(M1[31:30]));

wire [2:0] layer0_N16_wire = {M0[389], M0[388], M0[381]};
layer0_N16 layer0_N16_inst (.M0(layer0_N16_wire), .M1(M1[33:32]));

wire [2:0] layer0_N17_wire = {M0[486], M0[424], M0[150]};
layer0_N17 layer0_N17_inst (.M0(layer0_N17_wire), .M1(M1[35:34]));

wire [2:0] layer0_N18_wire = {M0[391], M0[266], M0[40]};
layer0_N18 layer0_N18_inst (.M0(layer0_N18_wire), .M1(M1[37:36]));

wire [2:0] layer0_N19_wire = {M0[506], M0[434], M0[247]};
layer0_N19 layer0_N19_inst (.M0(layer0_N19_wire), .M1(M1[39:38]));

wire [2:0] layer0_N20_wire = {M0[278], M0[206], M0[147]};
layer0_N20 layer0_N20_inst (.M0(layer0_N20_wire), .M1(M1[41:40]));

wire [2:0] layer0_N21_wire = {M0[456], M0[452], M0[168]};
layer0_N21 layer0_N21_inst (.M0(layer0_N21_wire), .M1(M1[43:42]));

wire [2:0] layer0_N22_wire = {M0[237], M0[230], M0[6]};
layer0_N22 layer0_N22_inst (.M0(layer0_N22_wire), .M1(M1[45:44]));

wire [2:0] layer0_N23_wire = {M0[146], M0[137], M0[80]};
layer0_N23 layer0_N23_inst (.M0(layer0_N23_wire), .M1(M1[47:46]));

wire [2:0] layer0_N24_wire = {M0[455], M0[342], M0[147]};
layer0_N24 layer0_N24_inst (.M0(layer0_N24_wire), .M1(M1[49:48]));

wire [2:0] layer0_N25_wire = {M0[451], M0[446], M0[48]};
layer0_N25 layer0_N25_inst (.M0(layer0_N25_wire), .M1(M1[51:50]));

wire [2:0] layer0_N26_wire = {M0[505], M0[172], M0[158]};
layer0_N26 layer0_N26_inst (.M0(layer0_N26_wire), .M1(M1[53:52]));

wire [2:0] layer0_N27_wire = {M0[245], M0[68], M0[47]};
layer0_N27 layer0_N27_inst (.M0(layer0_N27_wire), .M1(M1[55:54]));

wire [2:0] layer0_N28_wire = {M0[361], M0[345], M0[129]};
layer0_N28 layer0_N28_inst (.M0(layer0_N28_wire), .M1(M1[57:56]));

wire [2:0] layer0_N29_wire = {M0[490], M0[196], M0[117]};
layer0_N29 layer0_N29_inst (.M0(layer0_N29_wire), .M1(M1[59:58]));

wire [2:0] layer0_N30_wire = {M0[500], M0[450], M0[172]};
layer0_N30 layer0_N30_inst (.M0(layer0_N30_wire), .M1(M1[61:60]));

wire [2:0] layer0_N31_wire = {M0[435], M0[267], M0[52]};
layer0_N31 layer0_N31_inst (.M0(layer0_N31_wire), .M1(M1[63:62]));

wire [2:0] layer0_N32_wire = {M0[270], M0[242], M0[179]};
layer0_N32 layer0_N32_inst (.M0(layer0_N32_wire), .M1(M1[65:64]));

wire [2:0] layer0_N33_wire = {M0[467], M0[425], M0[134]};
layer0_N33 layer0_N33_inst (.M0(layer0_N33_wire), .M1(M1[67:66]));

wire [2:0] layer0_N34_wire = {M0[494], M0[402], M0[289]};
layer0_N34 layer0_N34_inst (.M0(layer0_N34_wire), .M1(M1[69:68]));

wire [2:0] layer0_N35_wire = {M0[503], M0[254], M0[57]};
layer0_N35 layer0_N35_inst (.M0(layer0_N35_wire), .M1(M1[71:70]));

wire [2:0] layer0_N36_wire = {M0[500], M0[306], M0[81]};
layer0_N36 layer0_N36_inst (.M0(layer0_N36_wire), .M1(M1[73:72]));

wire [2:0] layer0_N37_wire = {M0[416], M0[108], M0[81]};
layer0_N37 layer0_N37_inst (.M0(layer0_N37_wire), .M1(M1[75:74]));

wire [2:0] layer0_N38_wire = {M0[206], M0[130], M0[39]};
layer0_N38 layer0_N38_inst (.M0(layer0_N38_wire), .M1(M1[77:76]));

wire [2:0] layer0_N39_wire = {M0[500], M0[263], M0[32]};
layer0_N39 layer0_N39_inst (.M0(layer0_N39_wire), .M1(M1[79:78]));

wire [2:0] layer0_N40_wire = {M0[403], M0[332], M0[0]};
layer0_N40 layer0_N40_inst (.M0(layer0_N40_wire), .M1(M1[81:80]));

wire [2:0] layer0_N41_wire = {M0[326], M0[176], M0[20]};
layer0_N41 layer0_N41_inst (.M0(layer0_N41_wire), .M1(M1[83:82]));

wire [2:0] layer0_N42_wire = {M0[437], M0[395], M0[337]};
layer0_N42 layer0_N42_inst (.M0(layer0_N42_wire), .M1(M1[85:84]));

wire [2:0] layer0_N43_wire = {M0[306], M0[182], M0[33]};
layer0_N43 layer0_N43_inst (.M0(layer0_N43_wire), .M1(M1[87:86]));

wire [2:0] layer0_N44_wire = {M0[509], M0[371], M0[16]};
layer0_N44 layer0_N44_inst (.M0(layer0_N44_wire), .M1(M1[89:88]));

wire [2:0] layer0_N45_wire = {M0[207], M0[183], M0[32]};
layer0_N45 layer0_N45_inst (.M0(layer0_N45_wire), .M1(M1[91:90]));

wire [2:0] layer0_N46_wire = {M0[323], M0[306], M0[159]};
layer0_N46 layer0_N46_inst (.M0(layer0_N46_wire), .M1(M1[93:92]));

wire [2:0] layer0_N47_wire = {M0[490], M0[427], M0[122]};
layer0_N47 layer0_N47_inst (.M0(layer0_N47_wire), .M1(M1[95:94]));

wire [2:0] layer0_N48_wire = {M0[437], M0[248], M0[99]};
layer0_N48 layer0_N48_inst (.M0(layer0_N48_wire), .M1(M1[97:96]));

wire [2:0] layer0_N49_wire = {M0[362], M0[171], M0[54]};
layer0_N49 layer0_N49_inst (.M0(layer0_N49_wire), .M1(M1[99:98]));

wire [2:0] layer0_N50_wire = {M0[270], M0[263], M0[21]};
layer0_N50 layer0_N50_inst (.M0(layer0_N50_wire), .M1(M1[101:100]));

wire [2:0] layer0_N51_wire = {M0[304], M0[138], M0[131]};
layer0_N51 layer0_N51_inst (.M0(layer0_N51_wire), .M1(M1[103:102]));

wire [2:0] layer0_N52_wire = {M0[456], M0[240], M0[90]};
layer0_N52 layer0_N52_inst (.M0(layer0_N52_wire), .M1(M1[105:104]));

wire [2:0] layer0_N53_wire = {M0[433], M0[239], M0[169]};
layer0_N53 layer0_N53_inst (.M0(layer0_N53_wire), .M1(M1[107:106]));

wire [2:0] layer0_N54_wire = {M0[352], M0[98], M0[9]};
layer0_N54 layer0_N54_inst (.M0(layer0_N54_wire), .M1(M1[109:108]));

wire [2:0] layer0_N55_wire = {M0[328], M0[282], M0[57]};
layer0_N55 layer0_N55_inst (.M0(layer0_N55_wire), .M1(M1[111:110]));

wire [2:0] layer0_N56_wire = {M0[77], M0[67], M0[11]};
layer0_N56 layer0_N56_inst (.M0(layer0_N56_wire), .M1(M1[113:112]));

wire [2:0] layer0_N57_wire = {M0[407], M0[328], M0[275]};
layer0_N57 layer0_N57_inst (.M0(layer0_N57_wire), .M1(M1[115:114]));

wire [2:0] layer0_N58_wire = {M0[475], M0[441], M0[100]};
layer0_N58 layer0_N58_inst (.M0(layer0_N58_wire), .M1(M1[117:116]));

wire [2:0] layer0_N59_wire = {M0[424], M0[348], M0[170]};
layer0_N59 layer0_N59_inst (.M0(layer0_N59_wire), .M1(M1[119:118]));

wire [2:0] layer0_N60_wire = {M0[472], M0[288], M0[138]};
layer0_N60 layer0_N60_inst (.M0(layer0_N60_wire), .M1(M1[121:120]));

wire [2:0] layer0_N61_wire = {M0[232], M0[58], M0[3]};
layer0_N61 layer0_N61_inst (.M0(layer0_N61_wire), .M1(M1[123:122]));

wire [2:0] layer0_N62_wire = {M0[418], M0[383], M0[99]};
layer0_N62 layer0_N62_inst (.M0(layer0_N62_wire), .M1(M1[125:124]));

wire [2:0] layer0_N63_wire = {M0[447], M0[407], M0[150]};
layer0_N63 layer0_N63_inst (.M0(layer0_N63_wire), .M1(M1[127:126]));

wire [2:0] layer0_N64_wire = {M0[438], M0[370], M0[283]};
layer0_N64 layer0_N64_inst (.M0(layer0_N64_wire), .M1(M1[129:128]));

wire [2:0] layer0_N65_wire = {M0[317], M0[93], M0[80]};
layer0_N65 layer0_N65_inst (.M0(layer0_N65_wire), .M1(M1[131:130]));

wire [2:0] layer0_N66_wire = {M0[273], M0[250], M0[49]};
layer0_N66 layer0_N66_inst (.M0(layer0_N66_wire), .M1(M1[133:132]));

wire [2:0] layer0_N67_wire = {M0[492], M0[443], M0[208]};
layer0_N67 layer0_N67_inst (.M0(layer0_N67_wire), .M1(M1[135:134]));

wire [2:0] layer0_N68_wire = {M0[409], M0[279], M0[43]};
layer0_N68 layer0_N68_inst (.M0(layer0_N68_wire), .M1(M1[137:136]));

wire [2:0] layer0_N69_wire = {M0[449], M0[390], M0[83]};
layer0_N69 layer0_N69_inst (.M0(layer0_N69_wire), .M1(M1[139:138]));

wire [2:0] layer0_N70_wire = {M0[457], M0[218], M0[47]};
layer0_N70 layer0_N70_inst (.M0(layer0_N70_wire), .M1(M1[141:140]));

wire [2:0] layer0_N71_wire = {M0[355], M0[264], M0[216]};
layer0_N71 layer0_N71_inst (.M0(layer0_N71_wire), .M1(M1[143:142]));

wire [2:0] layer0_N72_wire = {M0[416], M0[209], M0[91]};
layer0_N72 layer0_N72_inst (.M0(layer0_N72_wire), .M1(M1[145:144]));

wire [2:0] layer0_N73_wire = {M0[345], M0[178], M0[32]};
layer0_N73 layer0_N73_inst (.M0(layer0_N73_wire), .M1(M1[147:146]));

wire [2:0] layer0_N74_wire = {M0[327], M0[293], M0[49]};
layer0_N74 layer0_N74_inst (.M0(layer0_N74_wire), .M1(M1[149:148]));

wire [2:0] layer0_N75_wire = {M0[422], M0[258], M0[93]};
layer0_N75 layer0_N75_inst (.M0(layer0_N75_wire), .M1(M1[151:150]));

wire [2:0] layer0_N76_wire = {M0[375], M0[347], M0[157]};
layer0_N76 layer0_N76_inst (.M0(layer0_N76_wire), .M1(M1[153:152]));

wire [2:0] layer0_N77_wire = {M0[425], M0[363], M0[202]};
layer0_N77 layer0_N77_inst (.M0(layer0_N77_wire), .M1(M1[155:154]));

wire [2:0] layer0_N78_wire = {M0[257], M0[176], M0[21]};
layer0_N78 layer0_N78_inst (.M0(layer0_N78_wire), .M1(M1[157:156]));

wire [2:0] layer0_N79_wire = {M0[234], M0[224], M0[156]};
layer0_N79 layer0_N79_inst (.M0(layer0_N79_wire), .M1(M1[159:158]));

wire [2:0] layer0_N80_wire = {M0[482], M0[371], M0[62]};
layer0_N80 layer0_N80_inst (.M0(layer0_N80_wire), .M1(M1[161:160]));

wire [2:0] layer0_N81_wire = {M0[456], M0[392], M0[38]};
layer0_N81 layer0_N81_inst (.M0(layer0_N81_wire), .M1(M1[163:162]));

wire [2:0] layer0_N82_wire = {M0[166], M0[157], M0[8]};
layer0_N82 layer0_N82_inst (.M0(layer0_N82_wire), .M1(M1[165:164]));

wire [2:0] layer0_N83_wire = {M0[468], M0[274], M0[217]};
layer0_N83 layer0_N83_inst (.M0(layer0_N83_wire), .M1(M1[167:166]));

wire [2:0] layer0_N84_wire = {M0[247], M0[116], M0[64]};
layer0_N84 layer0_N84_inst (.M0(layer0_N84_wire), .M1(M1[169:168]));

wire [2:0] layer0_N85_wire = {M0[382], M0[81], M0[51]};
layer0_N85 layer0_N85_inst (.M0(layer0_N85_wire), .M1(M1[171:170]));

wire [2:0] layer0_N86_wire = {M0[368], M0[343], M0[213]};
layer0_N86 layer0_N86_inst (.M0(layer0_N86_wire), .M1(M1[173:172]));

wire [2:0] layer0_N87_wire = {M0[435], M0[384], M0[24]};
layer0_N87 layer0_N87_inst (.M0(layer0_N87_wire), .M1(M1[175:174]));

wire [2:0] layer0_N88_wire = {M0[450], M0[270], M0[90]};
layer0_N88 layer0_N88_inst (.M0(layer0_N88_wire), .M1(M1[177:176]));

wire [2:0] layer0_N89_wire = {M0[496], M0[412], M0[134]};
layer0_N89 layer0_N89_inst (.M0(layer0_N89_wire), .M1(M1[179:178]));

wire [2:0] layer0_N90_wire = {M0[505], M0[197], M0[148]};
layer0_N90 layer0_N90_inst (.M0(layer0_N90_wire), .M1(M1[181:180]));

wire [2:0] layer0_N91_wire = {M0[462], M0[345], M0[319]};
layer0_N91 layer0_N91_inst (.M0(layer0_N91_wire), .M1(M1[183:182]));

wire [2:0] layer0_N92_wire = {M0[237], M0[186], M0[141]};
layer0_N92 layer0_N92_inst (.M0(layer0_N92_wire), .M1(M1[185:184]));

wire [2:0] layer0_N93_wire = {M0[436], M0[216], M0[173]};
layer0_N93 layer0_N93_inst (.M0(layer0_N93_wire), .M1(M1[187:186]));

wire [2:0] layer0_N94_wire = {M0[443], M0[397], M0[13]};
layer0_N94 layer0_N94_inst (.M0(layer0_N94_wire), .M1(M1[189:188]));

wire [2:0] layer0_N95_wire = {M0[284], M0[150], M0[54]};
layer0_N95 layer0_N95_inst (.M0(layer0_N95_wire), .M1(M1[191:190]));

wire [2:0] layer0_N96_wire = {M0[221], M0[44], M0[16]};
layer0_N96 layer0_N96_inst (.M0(layer0_N96_wire), .M1(M1[193:192]));

wire [2:0] layer0_N97_wire = {M0[469], M0[368], M0[85]};
layer0_N97 layer0_N97_inst (.M0(layer0_N97_wire), .M1(M1[195:194]));

wire [2:0] layer0_N98_wire = {M0[118], M0[35], M0[24]};
layer0_N98 layer0_N98_inst (.M0(layer0_N98_wire), .M1(M1[197:196]));

wire [2:0] layer0_N99_wire = {M0[510], M0[155], M0[64]};
layer0_N99 layer0_N99_inst (.M0(layer0_N99_wire), .M1(M1[199:198]));

wire [2:0] layer0_N100_wire = {M0[467], M0[289], M0[62]};
layer0_N100 layer0_N100_inst (.M0(layer0_N100_wire), .M1(M1[201:200]));

wire [2:0] layer0_N101_wire = {M0[440], M0[276], M0[17]};
layer0_N101 layer0_N101_inst (.M0(layer0_N101_wire), .M1(M1[203:202]));

wire [2:0] layer0_N102_wire = {M0[302], M0[237], M0[9]};
layer0_N102 layer0_N102_inst (.M0(layer0_N102_wire), .M1(M1[205:204]));

wire [2:0] layer0_N103_wire = {M0[460], M0[150], M0[19]};
layer0_N103 layer0_N103_inst (.M0(layer0_N103_wire), .M1(M1[207:206]));

wire [2:0] layer0_N104_wire = {M0[407], M0[341], M0[112]};
layer0_N104 layer0_N104_inst (.M0(layer0_N104_wire), .M1(M1[209:208]));

wire [2:0] layer0_N105_wire = {M0[334], M0[286], M0[192]};
layer0_N105 layer0_N105_inst (.M0(layer0_N105_wire), .M1(M1[211:210]));

wire [2:0] layer0_N106_wire = {M0[490], M0[296], M0[187]};
layer0_N106 layer0_N106_inst (.M0(layer0_N106_wire), .M1(M1[213:212]));

wire [2:0] layer0_N107_wire = {M0[320], M0[273], M0[162]};
layer0_N107 layer0_N107_inst (.M0(layer0_N107_wire), .M1(M1[215:214]));

wire [2:0] layer0_N108_wire = {M0[391], M0[142], M0[33]};
layer0_N108 layer0_N108_inst (.M0(layer0_N108_wire), .M1(M1[217:216]));

wire [2:0] layer0_N109_wire = {M0[470], M0[422], M0[410]};
layer0_N109 layer0_N109_inst (.M0(layer0_N109_wire), .M1(M1[219:218]));

wire [2:0] layer0_N110_wire = {M0[507], M0[218], M0[216]};
layer0_N110 layer0_N110_inst (.M0(layer0_N110_wire), .M1(M1[221:220]));

wire [2:0] layer0_N111_wire = {M0[208], M0[148], M0[2]};
layer0_N111 layer0_N111_inst (.M0(layer0_N111_wire), .M1(M1[223:222]));

wire [2:0] layer0_N112_wire = {M0[380], M0[217], M0[68]};
layer0_N112 layer0_N112_inst (.M0(layer0_N112_wire), .M1(M1[225:224]));

wire [2:0] layer0_N113_wire = {M0[469], M0[83], M0[4]};
layer0_N113 layer0_N113_inst (.M0(layer0_N113_wire), .M1(M1[227:226]));

wire [2:0] layer0_N114_wire = {M0[379], M0[310], M0[149]};
layer0_N114 layer0_N114_inst (.M0(layer0_N114_wire), .M1(M1[229:228]));

wire [2:0] layer0_N115_wire = {M0[399], M0[351], M0[98]};
layer0_N115 layer0_N115_inst (.M0(layer0_N115_wire), .M1(M1[231:230]));

wire [2:0] layer0_N116_wire = {M0[499], M0[403], M0[279]};
layer0_N116 layer0_N116_inst (.M0(layer0_N116_wire), .M1(M1[233:232]));

wire [2:0] layer0_N117_wire = {M0[504], M0[351], M0[206]};
layer0_N117 layer0_N117_inst (.M0(layer0_N117_wire), .M1(M1[235:234]));

wire [2:0] layer0_N118_wire = {M0[240], M0[205], M0[72]};
layer0_N118 layer0_N118_inst (.M0(layer0_N118_wire), .M1(M1[237:236]));

wire [2:0] layer0_N119_wire = {M0[354], M0[81], M0[71]};
layer0_N119 layer0_N119_inst (.M0(layer0_N119_wire), .M1(M1[239:238]));

wire [2:0] layer0_N120_wire = {M0[484], M0[160], M0[16]};
layer0_N120 layer0_N120_inst (.M0(layer0_N120_wire), .M1(M1[241:240]));

wire [2:0] layer0_N121_wire = {M0[446], M0[413], M0[311]};
layer0_N121 layer0_N121_inst (.M0(layer0_N121_wire), .M1(M1[243:242]));

wire [2:0] layer0_N122_wire = {M0[413], M0[258], M0[119]};
layer0_N122 layer0_N122_inst (.M0(layer0_N122_wire), .M1(M1[245:244]));

wire [2:0] layer0_N123_wire = {M0[314], M0[298], M0[29]};
layer0_N123 layer0_N123_inst (.M0(layer0_N123_wire), .M1(M1[247:246]));

wire [2:0] layer0_N124_wire = {M0[404], M0[392], M0[194]};
layer0_N124 layer0_N124_inst (.M0(layer0_N124_wire), .M1(M1[249:248]));

wire [2:0] layer0_N125_wire = {M0[463], M0[392], M0[43]};
layer0_N125 layer0_N125_inst (.M0(layer0_N125_wire), .M1(M1[251:250]));

wire [2:0] layer0_N126_wire = {M0[462], M0[461], M0[322]};
layer0_N126 layer0_N126_inst (.M0(layer0_N126_wire), .M1(M1[253:252]));

wire [2:0] layer0_N127_wire = {M0[444], M0[245], M0[15]};
layer0_N127 layer0_N127_inst (.M0(layer0_N127_wire), .M1(M1[255:254]));

wire [2:0] layer0_N128_wire = {M0[301], M0[249], M0[112]};
layer0_N128 layer0_N128_inst (.M0(layer0_N128_wire), .M1(M1[257:256]));

wire [2:0] layer0_N129_wire = {M0[360], M0[336], M0[327]};
layer0_N129 layer0_N129_inst (.M0(layer0_N129_wire), .M1(M1[259:258]));

wire [2:0] layer0_N130_wire = {M0[500], M0[358], M0[283]};
layer0_N130 layer0_N130_inst (.M0(layer0_N130_wire), .M1(M1[261:260]));

wire [2:0] layer0_N131_wire = {M0[501], M0[483], M0[231]};
layer0_N131 layer0_N131_inst (.M0(layer0_N131_wire), .M1(M1[263:262]));

wire [2:0] layer0_N132_wire = {M0[400], M0[165], M0[90]};
layer0_N132 layer0_N132_inst (.M0(layer0_N132_wire), .M1(M1[265:264]));

wire [2:0] layer0_N133_wire = {M0[287], M0[246], M0[59]};
layer0_N133 layer0_N133_inst (.M0(layer0_N133_wire), .M1(M1[267:266]));

wire [2:0] layer0_N134_wire = {M0[300], M0[171], M0[69]};
layer0_N134 layer0_N134_inst (.M0(layer0_N134_wire), .M1(M1[269:268]));

wire [2:0] layer0_N135_wire = {M0[511], M0[488], M0[239]};
layer0_N135 layer0_N135_inst (.M0(layer0_N135_wire), .M1(M1[271:270]));

wire [2:0] layer0_N136_wire = {M0[257], M0[188], M0[44]};
layer0_N136 layer0_N136_inst (.M0(layer0_N136_wire), .M1(M1[273:272]));

wire [2:0] layer0_N137_wire = {M0[221], M0[168], M0[94]};
layer0_N137 layer0_N137_inst (.M0(layer0_N137_wire), .M1(M1[275:274]));

wire [2:0] layer0_N138_wire = {M0[397], M0[319], M0[83]};
layer0_N138 layer0_N138_inst (.M0(layer0_N138_wire), .M1(M1[277:276]));

wire [2:0] layer0_N139_wire = {M0[480], M0[473], M0[238]};
layer0_N139 layer0_N139_inst (.M0(layer0_N139_wire), .M1(M1[279:278]));

wire [2:0] layer0_N140_wire = {M0[353], M0[299], M0[133]};
layer0_N140 layer0_N140_inst (.M0(layer0_N140_wire), .M1(M1[281:280]));

wire [2:0] layer0_N141_wire = {M0[492], M0[419], M0[353]};
layer0_N141 layer0_N141_inst (.M0(layer0_N141_wire), .M1(M1[283:282]));

wire [2:0] layer0_N142_wire = {M0[432], M0[236], M0[111]};
layer0_N142 layer0_N142_inst (.M0(layer0_N142_wire), .M1(M1[285:284]));

wire [2:0] layer0_N143_wire = {M0[285], M0[228], M0[41]};
layer0_N143 layer0_N143_inst (.M0(layer0_N143_wire), .M1(M1[287:286]));

wire [2:0] layer0_N144_wire = {M0[427], M0[404], M0[50]};
layer0_N144 layer0_N144_inst (.M0(layer0_N144_wire), .M1(M1[289:288]));

wire [2:0] layer0_N145_wire = {M0[425], M0[301], M0[130]};
layer0_N145 layer0_N145_inst (.M0(layer0_N145_wire), .M1(M1[291:290]));

wire [2:0] layer0_N146_wire = {M0[223], M0[200], M0[195]};
layer0_N146 layer0_N146_inst (.M0(layer0_N146_wire), .M1(M1[293:292]));

wire [2:0] layer0_N147_wire = {M0[462], M0[143], M0[65]};
layer0_N147 layer0_N147_inst (.M0(layer0_N147_wire), .M1(M1[295:294]));

wire [2:0] layer0_N148_wire = {M0[327], M0[164], M0[92]};
layer0_N148 layer0_N148_inst (.M0(layer0_N148_wire), .M1(M1[297:296]));

wire [2:0] layer0_N149_wire = {M0[450], M0[337], M0[334]};
layer0_N149 layer0_N149_inst (.M0(layer0_N149_wire), .M1(M1[299:298]));

wire [2:0] layer0_N150_wire = {M0[389], M0[322], M0[254]};
layer0_N150 layer0_N150_inst (.M0(layer0_N150_wire), .M1(M1[301:300]));

wire [2:0] layer0_N151_wire = {M0[407], M0[309], M0[244]};
layer0_N151 layer0_N151_inst (.M0(layer0_N151_wire), .M1(M1[303:302]));

wire [2:0] layer0_N152_wire = {M0[451], M0[347], M0[65]};
layer0_N152 layer0_N152_inst (.M0(layer0_N152_wire), .M1(M1[305:304]));

wire [2:0] layer0_N153_wire = {M0[482], M0[440], M0[316]};
layer0_N153 layer0_N153_inst (.M0(layer0_N153_wire), .M1(M1[307:306]));

wire [2:0] layer0_N154_wire = {M0[476], M0[326], M0[92]};
layer0_N154 layer0_N154_inst (.M0(layer0_N154_wire), .M1(M1[309:308]));

wire [2:0] layer0_N155_wire = {M0[461], M0[124], M0[26]};
layer0_N155 layer0_N155_inst (.M0(layer0_N155_wire), .M1(M1[311:310]));

wire [2:0] layer0_N156_wire = {M0[163], M0[161], M0[138]};
layer0_N156 layer0_N156_inst (.M0(layer0_N156_wire), .M1(M1[313:312]));

wire [2:0] layer0_N157_wire = {M0[19], M0[7], M0[5]};
layer0_N157 layer0_N157_inst (.M0(layer0_N157_wire), .M1(M1[315:314]));

wire [2:0] layer0_N158_wire = {M0[339], M0[87], M0[49]};
layer0_N158 layer0_N158_inst (.M0(layer0_N158_wire), .M1(M1[317:316]));

wire [2:0] layer0_N159_wire = {M0[436], M0[294], M0[77]};
layer0_N159 layer0_N159_inst (.M0(layer0_N159_wire), .M1(M1[319:318]));

wire [2:0] layer0_N160_wire = {M0[192], M0[129], M0[110]};
layer0_N160 layer0_N160_inst (.M0(layer0_N160_wire), .M1(M1[321:320]));

wire [2:0] layer0_N161_wire = {M0[369], M0[244], M0[101]};
layer0_N161 layer0_N161_inst (.M0(layer0_N161_wire), .M1(M1[323:322]));

wire [2:0] layer0_N162_wire = {M0[478], M0[435], M0[180]};
layer0_N162 layer0_N162_inst (.M0(layer0_N162_wire), .M1(M1[325:324]));

wire [2:0] layer0_N163_wire = {M0[384], M0[110], M0[78]};
layer0_N163 layer0_N163_inst (.M0(layer0_N163_wire), .M1(M1[327:326]));

wire [2:0] layer0_N164_wire = {M0[307], M0[265], M0[249]};
layer0_N164 layer0_N164_inst (.M0(layer0_N164_wire), .M1(M1[329:328]));

wire [2:0] layer0_N165_wire = {M0[495], M0[353], M0[257]};
layer0_N165 layer0_N165_inst (.M0(layer0_N165_wire), .M1(M1[331:330]));

wire [2:0] layer0_N166_wire = {M0[381], M0[182], M0[65]};
layer0_N166 layer0_N166_inst (.M0(layer0_N166_wire), .M1(M1[333:332]));

wire [2:0] layer0_N167_wire = {M0[208], M0[182], M0[142]};
layer0_N167 layer0_N167_inst (.M0(layer0_N167_wire), .M1(M1[335:334]));

wire [2:0] layer0_N168_wire = {M0[414], M0[291], M0[196]};
layer0_N168 layer0_N168_inst (.M0(layer0_N168_wire), .M1(M1[337:336]));

wire [2:0] layer0_N169_wire = {M0[316], M0[264], M0[150]};
layer0_N169 layer0_N169_inst (.M0(layer0_N169_wire), .M1(M1[339:338]));

wire [2:0] layer0_N170_wire = {M0[207], M0[101], M0[24]};
layer0_N170 layer0_N170_inst (.M0(layer0_N170_wire), .M1(M1[341:340]));

wire [2:0] layer0_N171_wire = {M0[294], M0[281], M0[86]};
layer0_N171 layer0_N171_inst (.M0(layer0_N171_wire), .M1(M1[343:342]));

wire [2:0] layer0_N172_wire = {M0[339], M0[168], M0[48]};
layer0_N172 layer0_N172_inst (.M0(layer0_N172_wire), .M1(M1[345:344]));

wire [2:0] layer0_N173_wire = {M0[464], M0[190], M0[73]};
layer0_N173 layer0_N173_inst (.M0(layer0_N173_wire), .M1(M1[347:346]));

wire [2:0] layer0_N174_wire = {M0[351], M0[325], M0[295]};
layer0_N174 layer0_N174_inst (.M0(layer0_N174_wire), .M1(M1[349:348]));

wire [2:0] layer0_N175_wire = {M0[233], M0[209], M0[23]};
layer0_N175 layer0_N175_inst (.M0(layer0_N175_wire), .M1(M1[351:350]));

wire [2:0] layer0_N176_wire = {M0[505], M0[241], M0[8]};
layer0_N176 layer0_N176_inst (.M0(layer0_N176_wire), .M1(M1[353:352]));

wire [2:0] layer0_N177_wire = {M0[436], M0[401], M0[380]};
layer0_N177 layer0_N177_inst (.M0(layer0_N177_wire), .M1(M1[355:354]));

wire [2:0] layer0_N178_wire = {M0[122], M0[54], M0[13]};
layer0_N178 layer0_N178_inst (.M0(layer0_N178_wire), .M1(M1[357:356]));

wire [2:0] layer0_N179_wire = {M0[488], M0[241], M0[214]};
layer0_N179 layer0_N179_inst (.M0(layer0_N179_wire), .M1(M1[359:358]));

wire [2:0] layer0_N180_wire = {M0[509], M0[447], M0[207]};
layer0_N180 layer0_N180_inst (.M0(layer0_N180_wire), .M1(M1[361:360]));

wire [2:0] layer0_N181_wire = {M0[177], M0[167], M0[165]};
layer0_N181 layer0_N181_inst (.M0(layer0_N181_wire), .M1(M1[363:362]));

wire [2:0] layer0_N182_wire = {M0[288], M0[138], M0[8]};
layer0_N182 layer0_N182_inst (.M0(layer0_N182_wire), .M1(M1[365:364]));

wire [2:0] layer0_N183_wire = {M0[474], M0[443], M0[349]};
layer0_N183 layer0_N183_inst (.M0(layer0_N183_wire), .M1(M1[367:366]));

wire [2:0] layer0_N184_wire = {M0[433], M0[268], M0[210]};
layer0_N184 layer0_N184_inst (.M0(layer0_N184_wire), .M1(M1[369:368]));

wire [2:0] layer0_N185_wire = {M0[328], M0[261], M0[15]};
layer0_N185 layer0_N185_inst (.M0(layer0_N185_wire), .M1(M1[371:370]));

wire [2:0] layer0_N186_wire = {M0[454], M0[304], M0[163]};
layer0_N186 layer0_N186_inst (.M0(layer0_N186_wire), .M1(M1[373:372]));

wire [2:0] layer0_N187_wire = {M0[500], M0[449], M0[76]};
layer0_N187 layer0_N187_inst (.M0(layer0_N187_wire), .M1(M1[375:374]));

wire [2:0] layer0_N188_wire = {M0[201], M0[27], M0[23]};
layer0_N188 layer0_N188_inst (.M0(layer0_N188_wire), .M1(M1[377:376]));

wire [2:0] layer0_N189_wire = {M0[282], M0[190], M0[146]};
layer0_N189 layer0_N189_inst (.M0(layer0_N189_wire), .M1(M1[379:378]));

wire [2:0] layer0_N190_wire = {M0[482], M0[435], M0[99]};
layer0_N190 layer0_N190_inst (.M0(layer0_N190_wire), .M1(M1[381:380]));

wire [2:0] layer0_N191_wire = {M0[487], M0[474], M0[300]};
layer0_N191 layer0_N191_inst (.M0(layer0_N191_wire), .M1(M1[383:382]));

wire [2:0] layer0_N192_wire = {M0[379], M0[342], M0[190]};
layer0_N192 layer0_N192_inst (.M0(layer0_N192_wire), .M1(M1[385:384]));

wire [2:0] layer0_N193_wire = {M0[452], M0[403], M0[308]};
layer0_N193 layer0_N193_inst (.M0(layer0_N193_wire), .M1(M1[387:386]));

wire [2:0] layer0_N194_wire = {M0[471], M0[362], M0[329]};
layer0_N194 layer0_N194_inst (.M0(layer0_N194_wire), .M1(M1[389:388]));

wire [2:0] layer0_N195_wire = {M0[487], M0[158], M0[145]};
layer0_N195 layer0_N195_inst (.M0(layer0_N195_wire), .M1(M1[391:390]));

wire [2:0] layer0_N196_wire = {M0[214], M0[174], M0[21]};
layer0_N196 layer0_N196_inst (.M0(layer0_N196_wire), .M1(M1[393:392]));

wire [2:0] layer0_N197_wire = {M0[364], M0[332], M0[58]};
layer0_N197 layer0_N197_inst (.M0(layer0_N197_wire), .M1(M1[395:394]));

wire [2:0] layer0_N198_wire = {M0[431], M0[386], M0[269]};
layer0_N198 layer0_N198_inst (.M0(layer0_N198_wire), .M1(M1[397:396]));

wire [2:0] layer0_N199_wire = {M0[496], M0[404], M0[351]};
layer0_N199 layer0_N199_inst (.M0(layer0_N199_wire), .M1(M1[399:398]));

wire [2:0] layer0_N200_wire = {M0[323], M0[110], M0[74]};
layer0_N200 layer0_N200_inst (.M0(layer0_N200_wire), .M1(M1[401:400]));

wire [2:0] layer0_N201_wire = {M0[317], M0[275], M0[63]};
layer0_N201 layer0_N201_inst (.M0(layer0_N201_wire), .M1(M1[403:402]));

wire [2:0] layer0_N202_wire = {M0[365], M0[226], M0[102]};
layer0_N202 layer0_N202_inst (.M0(layer0_N202_wire), .M1(M1[405:404]));

wire [2:0] layer0_N203_wire = {M0[393], M0[196], M0[50]};
layer0_N203 layer0_N203_inst (.M0(layer0_N203_wire), .M1(M1[407:406]));

wire [2:0] layer0_N204_wire = {M0[164], M0[118], M0[67]};
layer0_N204 layer0_N204_inst (.M0(layer0_N204_wire), .M1(M1[409:408]));

wire [2:0] layer0_N205_wire = {M0[496], M0[475], M0[463]};
layer0_N205 layer0_N205_inst (.M0(layer0_N205_wire), .M1(M1[411:410]));

wire [2:0] layer0_N206_wire = {M0[412], M0[268], M0[267]};
layer0_N206 layer0_N206_inst (.M0(layer0_N206_wire), .M1(M1[413:412]));

wire [2:0] layer0_N207_wire = {M0[309], M0[140], M0[123]};
layer0_N207 layer0_N207_inst (.M0(layer0_N207_wire), .M1(M1[415:414]));

wire [2:0] layer0_N208_wire = {M0[316], M0[53], M0[22]};
layer0_N208 layer0_N208_inst (.M0(layer0_N208_wire), .M1(M1[417:416]));

wire [2:0] layer0_N209_wire = {M0[385], M0[276], M0[130]};
layer0_N209 layer0_N209_inst (.M0(layer0_N209_wire), .M1(M1[419:418]));

wire [2:0] layer0_N210_wire = {M0[337], M0[327], M0[321]};
layer0_N210 layer0_N210_inst (.M0(layer0_N210_wire), .M1(M1[421:420]));

wire [2:0] layer0_N211_wire = {M0[459], M0[179], M0[150]};
layer0_N211 layer0_N211_inst (.M0(layer0_N211_wire), .M1(M1[423:422]));

wire [2:0] layer0_N212_wire = {M0[488], M0[350], M0[265]};
layer0_N212 layer0_N212_inst (.M0(layer0_N212_wire), .M1(M1[425:424]));

wire [2:0] layer0_N213_wire = {M0[364], M0[353], M0[199]};
layer0_N213 layer0_N213_inst (.M0(layer0_N213_wire), .M1(M1[427:426]));

wire [2:0] layer0_N214_wire = {M0[488], M0[289], M0[258]};
layer0_N214 layer0_N214_inst (.M0(layer0_N214_wire), .M1(M1[429:428]));

wire [2:0] layer0_N215_wire = {M0[484], M0[373], M0[355]};
layer0_N215 layer0_N215_inst (.M0(layer0_N215_wire), .M1(M1[431:430]));

wire [2:0] layer0_N216_wire = {M0[185], M0[64], M0[48]};
layer0_N216 layer0_N216_inst (.M0(layer0_N216_wire), .M1(M1[433:432]));

wire [2:0] layer0_N217_wire = {M0[78], M0[63], M0[31]};
layer0_N217 layer0_N217_inst (.M0(layer0_N217_wire), .M1(M1[435:434]));

wire [2:0] layer0_N218_wire = {M0[428], M0[418], M0[412]};
layer0_N218 layer0_N218_inst (.M0(layer0_N218_wire), .M1(M1[437:436]));

wire [2:0] layer0_N219_wire = {M0[491], M0[283], M0[176]};
layer0_N219 layer0_N219_inst (.M0(layer0_N219_wire), .M1(M1[439:438]));

wire [2:0] layer0_N220_wire = {M0[380], M0[184], M0[67]};
layer0_N220 layer0_N220_inst (.M0(layer0_N220_wire), .M1(M1[441:440]));

wire [2:0] layer0_N221_wire = {M0[475], M0[309], M0[144]};
layer0_N221 layer0_N221_inst (.M0(layer0_N221_wire), .M1(M1[443:442]));

wire [2:0] layer0_N222_wire = {M0[226], M0[65], M0[52]};
layer0_N222 layer0_N222_inst (.M0(layer0_N222_wire), .M1(M1[445:444]));

wire [2:0] layer0_N223_wire = {M0[398], M0[179], M0[41]};
layer0_N223 layer0_N223_inst (.M0(layer0_N223_wire), .M1(M1[447:446]));

wire [2:0] layer0_N224_wire = {M0[123], M0[49], M0[2]};
layer0_N224 layer0_N224_inst (.M0(layer0_N224_wire), .M1(M1[449:448]));

wire [2:0] layer0_N225_wire = {M0[371], M0[281], M0[47]};
layer0_N225 layer0_N225_inst (.M0(layer0_N225_wire), .M1(M1[451:450]));

wire [2:0] layer0_N226_wire = {M0[401], M0[369], M0[53]};
layer0_N226 layer0_N226_inst (.M0(layer0_N226_wire), .M1(M1[453:452]));

wire [2:0] layer0_N227_wire = {M0[486], M0[190], M0[48]};
layer0_N227 layer0_N227_inst (.M0(layer0_N227_wire), .M1(M1[455:454]));

wire [2:0] layer0_N228_wire = {M0[351], M0[11], M0[4]};
layer0_N228 layer0_N228_inst (.M0(layer0_N228_wire), .M1(M1[457:456]));

wire [2:0] layer0_N229_wire = {M0[493], M0[133], M0[120]};
layer0_N229 layer0_N229_inst (.M0(layer0_N229_wire), .M1(M1[459:458]));

wire [2:0] layer0_N230_wire = {M0[356], M0[237], M0[48]};
layer0_N230 layer0_N230_inst (.M0(layer0_N230_wire), .M1(M1[461:460]));

wire [2:0] layer0_N231_wire = {M0[199], M0[149], M0[20]};
layer0_N231 layer0_N231_inst (.M0(layer0_N231_wire), .M1(M1[463:462]));

wire [2:0] layer0_N232_wire = {M0[450], M0[346], M0[314]};
layer0_N232 layer0_N232_inst (.M0(layer0_N232_wire), .M1(M1[465:464]));

wire [2:0] layer0_N233_wire = {M0[503], M0[154], M0[23]};
layer0_N233 layer0_N233_inst (.M0(layer0_N233_wire), .M1(M1[467:466]));

wire [2:0] layer0_N234_wire = {M0[454], M0[341], M0[197]};
layer0_N234 layer0_N234_inst (.M0(layer0_N234_wire), .M1(M1[469:468]));

wire [2:0] layer0_N235_wire = {M0[313], M0[186], M0[56]};
layer0_N235 layer0_N235_inst (.M0(layer0_N235_wire), .M1(M1[471:470]));

wire [2:0] layer0_N236_wire = {M0[509], M0[375], M0[120]};
layer0_N236 layer0_N236_inst (.M0(layer0_N236_wire), .M1(M1[473:472]));

wire [2:0] layer0_N237_wire = {M0[296], M0[248], M0[61]};
layer0_N237 layer0_N237_inst (.M0(layer0_N237_wire), .M1(M1[475:474]));

wire [2:0] layer0_N238_wire = {M0[336], M0[310], M0[160]};
layer0_N238 layer0_N238_inst (.M0(layer0_N238_wire), .M1(M1[477:476]));

wire [2:0] layer0_N239_wire = {M0[471], M0[210], M0[102]};
layer0_N239 layer0_N239_inst (.M0(layer0_N239_wire), .M1(M1[479:478]));

wire [2:0] layer0_N240_wire = {M0[405], M0[341], M0[129]};
layer0_N240 layer0_N240_inst (.M0(layer0_N240_wire), .M1(M1[481:480]));

wire [2:0] layer0_N241_wire = {M0[317], M0[102], M0[70]};
layer0_N241 layer0_N241_inst (.M0(layer0_N241_wire), .M1(M1[483:482]));

wire [2:0] layer0_N242_wire = {M0[355], M0[306], M0[265]};
layer0_N242 layer0_N242_inst (.M0(layer0_N242_wire), .M1(M1[485:484]));

wire [2:0] layer0_N243_wire = {M0[434], M0[250], M0[1]};
layer0_N243 layer0_N243_inst (.M0(layer0_N243_wire), .M1(M1[487:486]));

wire [2:0] layer0_N244_wire = {M0[499], M0[355], M0[93]};
layer0_N244 layer0_N244_inst (.M0(layer0_N244_wire), .M1(M1[489:488]));

wire [2:0] layer0_N245_wire = {M0[406], M0[317], M0[121]};
layer0_N245 layer0_N245_inst (.M0(layer0_N245_wire), .M1(M1[491:490]));

wire [2:0] layer0_N246_wire = {M0[422], M0[73], M0[66]};
layer0_N246 layer0_N246_inst (.M0(layer0_N246_wire), .M1(M1[493:492]));

wire [2:0] layer0_N247_wire = {M0[424], M0[87], M0[39]};
layer0_N247 layer0_N247_inst (.M0(layer0_N247_wire), .M1(M1[495:494]));

wire [2:0] layer0_N248_wire = {M0[242], M0[156], M0[21]};
layer0_N248 layer0_N248_inst (.M0(layer0_N248_wire), .M1(M1[497:496]));

wire [2:0] layer0_N249_wire = {M0[498], M0[264], M0[51]};
layer0_N249 layer0_N249_inst (.M0(layer0_N249_wire), .M1(M1[499:498]));

wire [2:0] layer0_N250_wire = {M0[357], M0[162], M0[51]};
layer0_N250 layer0_N250_inst (.M0(layer0_N250_wire), .M1(M1[501:500]));

wire [2:0] layer0_N251_wire = {M0[403], M0[369], M0[311]};
layer0_N251 layer0_N251_inst (.M0(layer0_N251_wire), .M1(M1[503:502]));

wire [2:0] layer0_N252_wire = {M0[389], M0[155], M0[134]};
layer0_N252 layer0_N252_inst (.M0(layer0_N252_wire), .M1(M1[505:504]));

wire [2:0] layer0_N253_wire = {M0[485], M0[464], M0[140]};
layer0_N253 layer0_N253_inst (.M0(layer0_N253_wire), .M1(M1[507:506]));

wire [2:0] layer0_N254_wire = {M0[389], M0[195], M0[60]};
layer0_N254 layer0_N254_inst (.M0(layer0_N254_wire), .M1(M1[509:508]));

wire [2:0] layer0_N255_wire = {M0[464], M0[165], M0[128]};
layer0_N255 layer0_N255_inst (.M0(layer0_N255_wire), .M1(M1[511:510]));

wire [2:0] layer0_N256_wire = {M0[312], M0[262], M0[206]};
layer0_N256 layer0_N256_inst (.M0(layer0_N256_wire), .M1(M1[513:512]));

wire [2:0] layer0_N257_wire = {M0[441], M0[38], M0[3]};
layer0_N257 layer0_N257_inst (.M0(layer0_N257_wire), .M1(M1[515:514]));

wire [2:0] layer0_N258_wire = {M0[490], M0[147], M0[17]};
layer0_N258 layer0_N258_inst (.M0(layer0_N258_wire), .M1(M1[517:516]));

wire [2:0] layer0_N259_wire = {M0[107], M0[104], M0[62]};
layer0_N259 layer0_N259_inst (.M0(layer0_N259_wire), .M1(M1[519:518]));

wire [2:0] layer0_N260_wire = {M0[464], M0[448], M0[93]};
layer0_N260 layer0_N260_inst (.M0(layer0_N260_wire), .M1(M1[521:520]));

wire [2:0] layer0_N261_wire = {M0[391], M0[176], M0[39]};
layer0_N261 layer0_N261_inst (.M0(layer0_N261_wire), .M1(M1[523:522]));

wire [2:0] layer0_N262_wire = {M0[508], M0[104], M0[16]};
layer0_N262 layer0_N262_inst (.M0(layer0_N262_wire), .M1(M1[525:524]));

wire [2:0] layer0_N263_wire = {M0[441], M0[370], M0[266]};
layer0_N263 layer0_N263_inst (.M0(layer0_N263_wire), .M1(M1[527:526]));

wire [2:0] layer0_N264_wire = {M0[506], M0[473], M0[237]};
layer0_N264 layer0_N264_inst (.M0(layer0_N264_wire), .M1(M1[529:528]));

wire [2:0] layer0_N265_wire = {M0[459], M0[138], M0[131]};
layer0_N265 layer0_N265_inst (.M0(layer0_N265_wire), .M1(M1[531:530]));

wire [2:0] layer0_N266_wire = {M0[382], M0[297], M0[75]};
layer0_N266 layer0_N266_inst (.M0(layer0_N266_wire), .M1(M1[533:532]));

wire [2:0] layer0_N267_wire = {M0[353], M0[288], M0[234]};
layer0_N267 layer0_N267_inst (.M0(layer0_N267_wire), .M1(M1[535:534]));

wire [2:0] layer0_N268_wire = {M0[476], M0[212], M0[176]};
layer0_N268 layer0_N268_inst (.M0(layer0_N268_wire), .M1(M1[537:536]));

wire [2:0] layer0_N269_wire = {M0[474], M0[257], M0[62]};
layer0_N269 layer0_N269_inst (.M0(layer0_N269_wire), .M1(M1[539:538]));

wire [2:0] layer0_N270_wire = {M0[410], M0[220], M0[66]};
layer0_N270 layer0_N270_inst (.M0(layer0_N270_wire), .M1(M1[541:540]));

wire [2:0] layer0_N271_wire = {M0[112], M0[103], M0[79]};
layer0_N271 layer0_N271_inst (.M0(layer0_N271_wire), .M1(M1[543:542]));

wire [2:0] layer0_N272_wire = {M0[466], M0[374], M0[187]};
layer0_N272 layer0_N272_inst (.M0(layer0_N272_wire), .M1(M1[545:544]));

wire [2:0] layer0_N273_wire = {M0[495], M0[394], M0[278]};
layer0_N273 layer0_N273_inst (.M0(layer0_N273_wire), .M1(M1[547:546]));

wire [2:0] layer0_N274_wire = {M0[498], M0[151], M0[9]};
layer0_N274 layer0_N274_inst (.M0(layer0_N274_wire), .M1(M1[549:548]));

wire [2:0] layer0_N275_wire = {M0[335], M0[203], M0[29]};
layer0_N275 layer0_N275_inst (.M0(layer0_N275_wire), .M1(M1[551:550]));

wire [2:0] layer0_N276_wire = {M0[447], M0[285], M0[62]};
layer0_N276 layer0_N276_inst (.M0(layer0_N276_wire), .M1(M1[553:552]));

wire [2:0] layer0_N277_wire = {M0[353], M0[206], M0[34]};
layer0_N277 layer0_N277_inst (.M0(layer0_N277_wire), .M1(M1[555:554]));

wire [2:0] layer0_N278_wire = {M0[414], M0[347], M0[338]};
layer0_N278 layer0_N278_inst (.M0(layer0_N278_wire), .M1(M1[557:556]));

wire [2:0] layer0_N279_wire = {M0[261], M0[27], M0[23]};
layer0_N279 layer0_N279_inst (.M0(layer0_N279_wire), .M1(M1[559:558]));

wire [2:0] layer0_N280_wire = {M0[156], M0[151], M0[23]};
layer0_N280 layer0_N280_inst (.M0(layer0_N280_wire), .M1(M1[561:560]));

wire [2:0] layer0_N281_wire = {M0[337], M0[275], M0[97]};
layer0_N281 layer0_N281_inst (.M0(layer0_N281_wire), .M1(M1[563:562]));

wire [2:0] layer0_N282_wire = {M0[424], M0[325], M0[133]};
layer0_N282 layer0_N282_inst (.M0(layer0_N282_wire), .M1(M1[565:564]));

wire [2:0] layer0_N283_wire = {M0[497], M0[189], M0[125]};
layer0_N283 layer0_N283_inst (.M0(layer0_N283_wire), .M1(M1[567:566]));

wire [2:0] layer0_N284_wire = {M0[343], M0[192], M0[26]};
layer0_N284 layer0_N284_inst (.M0(layer0_N284_wire), .M1(M1[569:568]));

wire [2:0] layer0_N285_wire = {M0[402], M0[329], M0[269]};
layer0_N285 layer0_N285_inst (.M0(layer0_N285_wire), .M1(M1[571:570]));

wire [2:0] layer0_N286_wire = {M0[258], M0[254], M0[227]};
layer0_N286 layer0_N286_inst (.M0(layer0_N286_wire), .M1(M1[573:572]));

wire [2:0] layer0_N287_wire = {M0[312], M0[244], M0[147]};
layer0_N287 layer0_N287_inst (.M0(layer0_N287_wire), .M1(M1[575:574]));

wire [2:0] layer0_N288_wire = {M0[331], M0[305], M0[242]};
layer0_N288 layer0_N288_inst (.M0(layer0_N288_wire), .M1(M1[577:576]));

wire [2:0] layer0_N289_wire = {M0[509], M0[358], M0[348]};
layer0_N289 layer0_N289_inst (.M0(layer0_N289_wire), .M1(M1[579:578]));

wire [2:0] layer0_N290_wire = {M0[432], M0[402], M0[343]};
layer0_N290 layer0_N290_inst (.M0(layer0_N290_wire), .M1(M1[581:580]));

wire [2:0] layer0_N291_wire = {M0[499], M0[297], M0[255]};
layer0_N291 layer0_N291_inst (.M0(layer0_N291_wire), .M1(M1[583:582]));

wire [2:0] layer0_N292_wire = {M0[225], M0[154], M0[17]};
layer0_N292 layer0_N292_inst (.M0(layer0_N292_wire), .M1(M1[585:584]));

wire [2:0] layer0_N293_wire = {M0[401], M0[291], M0[268]};
layer0_N293 layer0_N293_inst (.M0(layer0_N293_wire), .M1(M1[587:586]));

wire [2:0] layer0_N294_wire = {M0[349], M0[323], M0[139]};
layer0_N294 layer0_N294_inst (.M0(layer0_N294_wire), .M1(M1[589:588]));

wire [2:0] layer0_N295_wire = {M0[400], M0[392], M0[276]};
layer0_N295 layer0_N295_inst (.M0(layer0_N295_wire), .M1(M1[591:590]));

wire [2:0] layer0_N296_wire = {M0[495], M0[394], M0[303]};
layer0_N296 layer0_N296_inst (.M0(layer0_N296_wire), .M1(M1[593:592]));

wire [2:0] layer0_N297_wire = {M0[449], M0[124], M0[91]};
layer0_N297 layer0_N297_inst (.M0(layer0_N297_wire), .M1(M1[595:594]));

wire [2:0] layer0_N298_wire = {M0[414], M0[211], M0[72]};
layer0_N298 layer0_N298_inst (.M0(layer0_N298_wire), .M1(M1[597:596]));

wire [2:0] layer0_N299_wire = {M0[195], M0[98], M0[4]};
layer0_N299 layer0_N299_inst (.M0(layer0_N299_wire), .M1(M1[599:598]));

wire [2:0] layer0_N300_wire = {M0[471], M0[68], M0[53]};
layer0_N300 layer0_N300_inst (.M0(layer0_N300_wire), .M1(M1[601:600]));

wire [2:0] layer0_N301_wire = {M0[490], M0[264], M0[231]};
layer0_N301 layer0_N301_inst (.M0(layer0_N301_wire), .M1(M1[603:602]));

wire [2:0] layer0_N302_wire = {M0[484], M0[470], M0[406]};
layer0_N302 layer0_N302_inst (.M0(layer0_N302_wire), .M1(M1[605:604]));

wire [2:0] layer0_N303_wire = {M0[309], M0[228], M0[84]};
layer0_N303 layer0_N303_inst (.M0(layer0_N303_wire), .M1(M1[607:606]));

wire [2:0] layer0_N304_wire = {M0[448], M0[415], M0[264]};
layer0_N304 layer0_N304_inst (.M0(layer0_N304_wire), .M1(M1[609:608]));

wire [2:0] layer0_N305_wire = {M0[432], M0[224], M0[48]};
layer0_N305 layer0_N305_inst (.M0(layer0_N305_wire), .M1(M1[611:610]));

wire [2:0] layer0_N306_wire = {M0[271], M0[261], M0[242]};
layer0_N306 layer0_N306_inst (.M0(layer0_N306_wire), .M1(M1[613:612]));

wire [2:0] layer0_N307_wire = {M0[503], M0[393], M0[383]};
layer0_N307 layer0_N307_inst (.M0(layer0_N307_wire), .M1(M1[615:614]));

wire [2:0] layer0_N308_wire = {M0[286], M0[178], M0[11]};
layer0_N308 layer0_N308_inst (.M0(layer0_N308_wire), .M1(M1[617:616]));

wire [2:0] layer0_N309_wire = {M0[186], M0[159], M0[76]};
layer0_N309 layer0_N309_inst (.M0(layer0_N309_wire), .M1(M1[619:618]));

wire [2:0] layer0_N310_wire = {M0[405], M0[343], M0[125]};
layer0_N310 layer0_N310_inst (.M0(layer0_N310_wire), .M1(M1[621:620]));

wire [2:0] layer0_N311_wire = {M0[458], M0[300], M0[283]};
layer0_N311 layer0_N311_inst (.M0(layer0_N311_wire), .M1(M1[623:622]));

wire [2:0] layer0_N312_wire = {M0[316], M0[244], M0[112]};
layer0_N312 layer0_N312_inst (.M0(layer0_N312_wire), .M1(M1[625:624]));

wire [2:0] layer0_N313_wire = {M0[427], M0[134], M0[74]};
layer0_N313 layer0_N313_inst (.M0(layer0_N313_wire), .M1(M1[627:626]));

wire [2:0] layer0_N314_wire = {M0[494], M0[90], M0[12]};
layer0_N314 layer0_N314_inst (.M0(layer0_N314_wire), .M1(M1[629:628]));

wire [2:0] layer0_N315_wire = {M0[434], M0[220], M0[101]};
layer0_N315 layer0_N315_inst (.M0(layer0_N315_wire), .M1(M1[631:630]));

wire [2:0] layer0_N316_wire = {M0[369], M0[164], M0[96]};
layer0_N316 layer0_N316_inst (.M0(layer0_N316_wire), .M1(M1[633:632]));

wire [2:0] layer0_N317_wire = {M0[373], M0[296], M0[178]};
layer0_N317 layer0_N317_inst (.M0(layer0_N317_wire), .M1(M1[635:634]));

wire [2:0] layer0_N318_wire = {M0[473], M0[179], M0[14]};
layer0_N318 layer0_N318_inst (.M0(layer0_N318_wire), .M1(M1[637:636]));

wire [2:0] layer0_N319_wire = {M0[367], M0[237], M0[232]};
layer0_N319 layer0_N319_inst (.M0(layer0_N319_wire), .M1(M1[639:638]));

wire [2:0] layer0_N320_wire = {M0[377], M0[128], M0[46]};
layer0_N320 layer0_N320_inst (.M0(layer0_N320_wire), .M1(M1[641:640]));

wire [2:0] layer0_N321_wire = {M0[357], M0[258], M0[198]};
layer0_N321 layer0_N321_inst (.M0(layer0_N321_wire), .M1(M1[643:642]));

wire [2:0] layer0_N322_wire = {M0[241], M0[118], M0[54]};
layer0_N322 layer0_N322_inst (.M0(layer0_N322_wire), .M1(M1[645:644]));

wire [2:0] layer0_N323_wire = {M0[443], M0[240], M0[19]};
layer0_N323 layer0_N323_inst (.M0(layer0_N323_wire), .M1(M1[647:646]));

wire [2:0] layer0_N324_wire = {M0[487], M0[396], M0[311]};
layer0_N324 layer0_N324_inst (.M0(layer0_N324_wire), .M1(M1[649:648]));

wire [2:0] layer0_N325_wire = {M0[282], M0[132], M0[48]};
layer0_N325 layer0_N325_inst (.M0(layer0_N325_wire), .M1(M1[651:650]));

wire [2:0] layer0_N326_wire = {M0[306], M0[184], M0[89]};
layer0_N326 layer0_N326_inst (.M0(layer0_N326_wire), .M1(M1[653:652]));

wire [2:0] layer0_N327_wire = {M0[427], M0[368], M0[261]};
layer0_N327 layer0_N327_inst (.M0(layer0_N327_wire), .M1(M1[655:654]));

wire [2:0] layer0_N328_wire = {M0[498], M0[324], M0[292]};
layer0_N328 layer0_N328_inst (.M0(layer0_N328_wire), .M1(M1[657:656]));

wire [2:0] layer0_N329_wire = {M0[239], M0[143], M0[13]};
layer0_N329 layer0_N329_inst (.M0(layer0_N329_wire), .M1(M1[659:658]));

wire [2:0] layer0_N330_wire = {M0[504], M0[456], M0[375]};
layer0_N330 layer0_N330_inst (.M0(layer0_N330_wire), .M1(M1[661:660]));

wire [2:0] layer0_N331_wire = {M0[284], M0[253], M0[75]};
layer0_N331 layer0_N331_inst (.M0(layer0_N331_wire), .M1(M1[663:662]));

wire [2:0] layer0_N332_wire = {M0[326], M0[257], M0[83]};
layer0_N332 layer0_N332_inst (.M0(layer0_N332_wire), .M1(M1[665:664]));

wire [2:0] layer0_N333_wire = {M0[498], M0[378], M0[55]};
layer0_N333 layer0_N333_inst (.M0(layer0_N333_wire), .M1(M1[667:666]));

wire [2:0] layer0_N334_wire = {M0[442], M0[262], M0[50]};
layer0_N334 layer0_N334_inst (.M0(layer0_N334_wire), .M1(M1[669:668]));

wire [2:0] layer0_N335_wire = {M0[260], M0[244], M0[66]};
layer0_N335 layer0_N335_inst (.M0(layer0_N335_wire), .M1(M1[671:670]));

wire [2:0] layer0_N336_wire = {M0[264], M0[251], M0[178]};
layer0_N336 layer0_N336_inst (.M0(layer0_N336_wire), .M1(M1[673:672]));

wire [2:0] layer0_N337_wire = {M0[271], M0[258], M0[165]};
layer0_N337 layer0_N337_inst (.M0(layer0_N337_wire), .M1(M1[675:674]));

wire [2:0] layer0_N338_wire = {M0[317], M0[314], M0[14]};
layer0_N338 layer0_N338_inst (.M0(layer0_N338_wire), .M1(M1[677:676]));

wire [2:0] layer0_N339_wire = {M0[360], M0[314], M0[312]};
layer0_N339 layer0_N339_inst (.M0(layer0_N339_wire), .M1(M1[679:678]));

wire [2:0] layer0_N340_wire = {M0[495], M0[474], M0[217]};
layer0_N340 layer0_N340_inst (.M0(layer0_N340_wire), .M1(M1[681:680]));

wire [2:0] layer0_N341_wire = {M0[405], M0[287], M0[96]};
layer0_N341 layer0_N341_inst (.M0(layer0_N341_wire), .M1(M1[683:682]));

wire [2:0] layer0_N342_wire = {M0[341], M0[251], M0[86]};
layer0_N342 layer0_N342_inst (.M0(layer0_N342_wire), .M1(M1[685:684]));

wire [2:0] layer0_N343_wire = {M0[301], M0[300], M0[39]};
layer0_N343 layer0_N343_inst (.M0(layer0_N343_wire), .M1(M1[687:686]));

wire [2:0] layer0_N344_wire = {M0[506], M0[119], M0[33]};
layer0_N344 layer0_N344_inst (.M0(layer0_N344_wire), .M1(M1[689:688]));

wire [2:0] layer0_N345_wire = {M0[501], M0[387], M0[273]};
layer0_N345 layer0_N345_inst (.M0(layer0_N345_wire), .M1(M1[691:690]));

wire [2:0] layer0_N346_wire = {M0[360], M0[81], M0[4]};
layer0_N346 layer0_N346_inst (.M0(layer0_N346_wire), .M1(M1[693:692]));

wire [2:0] layer0_N347_wire = {M0[303], M0[272], M0[254]};
layer0_N347 layer0_N347_inst (.M0(layer0_N347_wire), .M1(M1[695:694]));

wire [2:0] layer0_N348_wire = {M0[404], M0[180], M0[20]};
layer0_N348 layer0_N348_inst (.M0(layer0_N348_wire), .M1(M1[697:696]));

wire [2:0] layer0_N349_wire = {M0[279], M0[221], M0[72]};
layer0_N349 layer0_N349_inst (.M0(layer0_N349_wire), .M1(M1[699:698]));

wire [2:0] layer0_N350_wire = {M0[479], M0[399], M0[133]};
layer0_N350 layer0_N350_inst (.M0(layer0_N350_wire), .M1(M1[701:700]));

wire [2:0] layer0_N351_wire = {M0[414], M0[50], M0[47]};
layer0_N351 layer0_N351_inst (.M0(layer0_N351_wire), .M1(M1[703:702]));

wire [2:0] layer0_N352_wire = {M0[510], M0[460], M0[321]};
layer0_N352 layer0_N352_inst (.M0(layer0_N352_wire), .M1(M1[705:704]));

wire [2:0] layer0_N353_wire = {M0[377], M0[278], M0[32]};
layer0_N353 layer0_N353_inst (.M0(layer0_N353_wire), .M1(M1[707:706]));

wire [2:0] layer0_N354_wire = {M0[299], M0[209], M0[99]};
layer0_N354 layer0_N354_inst (.M0(layer0_N354_wire), .M1(M1[709:708]));

wire [2:0] layer0_N355_wire = {M0[231], M0[131], M0[51]};
layer0_N355 layer0_N355_inst (.M0(layer0_N355_wire), .M1(M1[711:710]));

wire [2:0] layer0_N356_wire = {M0[397], M0[359], M0[174]};
layer0_N356 layer0_N356_inst (.M0(layer0_N356_wire), .M1(M1[713:712]));

wire [2:0] layer0_N357_wire = {M0[483], M0[357], M0[96]};
layer0_N357 layer0_N357_inst (.M0(layer0_N357_wire), .M1(M1[715:714]));

wire [2:0] layer0_N358_wire = {M0[456], M0[307], M0[58]};
layer0_N358 layer0_N358_inst (.M0(layer0_N358_wire), .M1(M1[717:716]));

wire [2:0] layer0_N359_wire = {M0[300], M0[215], M0[120]};
layer0_N359 layer0_N359_inst (.M0(layer0_N359_wire), .M1(M1[719:718]));

wire [2:0] layer0_N360_wire = {M0[301], M0[72], M0[58]};
layer0_N360 layer0_N360_inst (.M0(layer0_N360_wire), .M1(M1[721:720]));

wire [2:0] layer0_N361_wire = {M0[396], M0[139], M0[15]};
layer0_N361 layer0_N361_inst (.M0(layer0_N361_wire), .M1(M1[723:722]));

wire [2:0] layer0_N362_wire = {M0[385], M0[351], M0[232]};
layer0_N362 layer0_N362_inst (.M0(layer0_N362_wire), .M1(M1[725:724]));

wire [2:0] layer0_N363_wire = {M0[505], M0[82], M0[47]};
layer0_N363 layer0_N363_inst (.M0(layer0_N363_wire), .M1(M1[727:726]));

wire [2:0] layer0_N364_wire = {M0[253], M0[208], M0[201]};
layer0_N364 layer0_N364_inst (.M0(layer0_N364_wire), .M1(M1[729:728]));

wire [2:0] layer0_N365_wire = {M0[492], M0[297], M0[188]};
layer0_N365 layer0_N365_inst (.M0(layer0_N365_wire), .M1(M1[731:730]));

wire [2:0] layer0_N366_wire = {M0[437], M0[358], M0[321]};
layer0_N366 layer0_N366_inst (.M0(layer0_N366_wire), .M1(M1[733:732]));

wire [2:0] layer0_N367_wire = {M0[216], M0[121], M0[112]};
layer0_N367 layer0_N367_inst (.M0(layer0_N367_wire), .M1(M1[735:734]));

wire [2:0] layer0_N368_wire = {M0[213], M0[61], M0[11]};
layer0_N368 layer0_N368_inst (.M0(layer0_N368_wire), .M1(M1[737:736]));

wire [2:0] layer0_N369_wire = {M0[403], M0[266], M0[188]};
layer0_N369 layer0_N369_inst (.M0(layer0_N369_wire), .M1(M1[739:738]));

wire [2:0] layer0_N370_wire = {M0[483], M0[143], M0[85]};
layer0_N370 layer0_N370_inst (.M0(layer0_N370_wire), .M1(M1[741:740]));

wire [2:0] layer0_N371_wire = {M0[495], M0[353], M0[245]};
layer0_N371 layer0_N371_inst (.M0(layer0_N371_wire), .M1(M1[743:742]));

wire [2:0] layer0_N372_wire = {M0[395], M0[297], M0[129]};
layer0_N372 layer0_N372_inst (.M0(layer0_N372_wire), .M1(M1[745:744]));

wire [2:0] layer0_N373_wire = {M0[491], M0[456], M0[9]};
layer0_N373 layer0_N373_inst (.M0(layer0_N373_wire), .M1(M1[747:746]));

wire [2:0] layer0_N374_wire = {M0[500], M0[199], M0[17]};
layer0_N374 layer0_N374_inst (.M0(layer0_N374_wire), .M1(M1[749:748]));

wire [2:0] layer0_N375_wire = {M0[256], M0[171], M0[161]};
layer0_N375 layer0_N375_inst (.M0(layer0_N375_wire), .M1(M1[751:750]));

wire [2:0] layer0_N376_wire = {M0[472], M0[384], M0[170]};
layer0_N376 layer0_N376_inst (.M0(layer0_N376_wire), .M1(M1[753:752]));

wire [2:0] layer0_N377_wire = {M0[229], M0[207], M0[178]};
layer0_N377 layer0_N377_inst (.M0(layer0_N377_wire), .M1(M1[755:754]));

wire [2:0] layer0_N378_wire = {M0[471], M0[86], M0[35]};
layer0_N378 layer0_N378_inst (.M0(layer0_N378_wire), .M1(M1[757:756]));

wire [2:0] layer0_N379_wire = {M0[316], M0[247], M0[165]};
layer0_N379 layer0_N379_inst (.M0(layer0_N379_wire), .M1(M1[759:758]));

wire [2:0] layer0_N380_wire = {M0[370], M0[351], M0[217]};
layer0_N380 layer0_N380_inst (.M0(layer0_N380_wire), .M1(M1[761:760]));

wire [2:0] layer0_N381_wire = {M0[357], M0[306], M0[162]};
layer0_N381 layer0_N381_inst (.M0(layer0_N381_wire), .M1(M1[763:762]));

wire [2:0] layer0_N382_wire = {M0[302], M0[163], M0[5]};
layer0_N382 layer0_N382_inst (.M0(layer0_N382_wire), .M1(M1[765:764]));

wire [2:0] layer0_N383_wire = {M0[475], M0[429], M0[351]};
layer0_N383 layer0_N383_inst (.M0(layer0_N383_wire), .M1(M1[767:766]));

wire [2:0] layer0_N384_wire = {M0[499], M0[428], M0[246]};
layer0_N384 layer0_N384_inst (.M0(layer0_N384_wire), .M1(M1[769:768]));

wire [2:0] layer0_N385_wire = {M0[347], M0[135], M0[127]};
layer0_N385 layer0_N385_inst (.M0(layer0_N385_wire), .M1(M1[771:770]));

wire [2:0] layer0_N386_wire = {M0[504], M0[248], M0[202]};
layer0_N386 layer0_N386_inst (.M0(layer0_N386_wire), .M1(M1[773:772]));

wire [2:0] layer0_N387_wire = {M0[450], M0[412], M0[20]};
layer0_N387 layer0_N387_inst (.M0(layer0_N387_wire), .M1(M1[775:774]));

wire [2:0] layer0_N388_wire = {M0[451], M0[315], M0[7]};
layer0_N388 layer0_N388_inst (.M0(layer0_N388_wire), .M1(M1[777:776]));

wire [2:0] layer0_N389_wire = {M0[298], M0[260], M0[128]};
layer0_N389 layer0_N389_inst (.M0(layer0_N389_wire), .M1(M1[779:778]));

wire [2:0] layer0_N390_wire = {M0[426], M0[375], M0[112]};
layer0_N390 layer0_N390_inst (.M0(layer0_N390_wire), .M1(M1[781:780]));

wire [2:0] layer0_N391_wire = {M0[379], M0[362], M0[146]};
layer0_N391 layer0_N391_inst (.M0(layer0_N391_wire), .M1(M1[783:782]));

wire [2:0] layer0_N392_wire = {M0[424], M0[190], M0[62]};
layer0_N392 layer0_N392_inst (.M0(layer0_N392_wire), .M1(M1[785:784]));

wire [2:0] layer0_N393_wire = {M0[491], M0[440], M0[199]};
layer0_N393 layer0_N393_inst (.M0(layer0_N393_wire), .M1(M1[787:786]));

wire [2:0] layer0_N394_wire = {M0[486], M0[125], M0[107]};
layer0_N394 layer0_N394_inst (.M0(layer0_N394_wire), .M1(M1[789:788]));

wire [2:0] layer0_N395_wire = {M0[277], M0[80], M0[56]};
layer0_N395 layer0_N395_inst (.M0(layer0_N395_wire), .M1(M1[791:790]));

wire [2:0] layer0_N396_wire = {M0[477], M0[369], M0[195]};
layer0_N396 layer0_N396_inst (.M0(layer0_N396_wire), .M1(M1[793:792]));

wire [2:0] layer0_N397_wire = {M0[475], M0[159], M0[9]};
layer0_N397 layer0_N397_inst (.M0(layer0_N397_wire), .M1(M1[795:794]));

wire [2:0] layer0_N398_wire = {M0[179], M0[72], M0[50]};
layer0_N398 layer0_N398_inst (.M0(layer0_N398_wire), .M1(M1[797:796]));

wire [2:0] layer0_N399_wire = {M0[475], M0[428], M0[45]};
layer0_N399 layer0_N399_inst (.M0(layer0_N399_wire), .M1(M1[799:798]));

wire [2:0] layer0_N400_wire = {M0[225], M0[60], M0[52]};
layer0_N400 layer0_N400_inst (.M0(layer0_N400_wire), .M1(M1[801:800]));

wire [2:0] layer0_N401_wire = {M0[458], M0[182], M0[103]};
layer0_N401 layer0_N401_inst (.M0(layer0_N401_wire), .M1(M1[803:802]));

wire [2:0] layer0_N402_wire = {M0[495], M0[466], M0[314]};
layer0_N402 layer0_N402_inst (.M0(layer0_N402_wire), .M1(M1[805:804]));

wire [2:0] layer0_N403_wire = {M0[498], M0[185], M0[82]};
layer0_N403 layer0_N403_inst (.M0(layer0_N403_wire), .M1(M1[807:806]));

wire [2:0] layer0_N404_wire = {M0[452], M0[361], M0[277]};
layer0_N404 layer0_N404_inst (.M0(layer0_N404_wire), .M1(M1[809:808]));

wire [2:0] layer0_N405_wire = {M0[240], M0[78], M0[24]};
layer0_N405 layer0_N405_inst (.M0(layer0_N405_wire), .M1(M1[811:810]));

wire [2:0] layer0_N406_wire = {M0[310], M0[257], M0[160]};
layer0_N406 layer0_N406_inst (.M0(layer0_N406_wire), .M1(M1[813:812]));

wire [2:0] layer0_N407_wire = {M0[410], M0[401], M0[303]};
layer0_N407 layer0_N407_inst (.M0(layer0_N407_wire), .M1(M1[815:814]));

wire [2:0] layer0_N408_wire = {M0[355], M0[221], M0[102]};
layer0_N408 layer0_N408_inst (.M0(layer0_N408_wire), .M1(M1[817:816]));

wire [2:0] layer0_N409_wire = {M0[342], M0[249], M0[131]};
layer0_N409 layer0_N409_inst (.M0(layer0_N409_wire), .M1(M1[819:818]));

wire [2:0] layer0_N410_wire = {M0[452], M0[397], M0[88]};
layer0_N410 layer0_N410_inst (.M0(layer0_N410_wire), .M1(M1[821:820]));

wire [2:0] layer0_N411_wire = {M0[371], M0[186], M0[25]};
layer0_N411 layer0_N411_inst (.M0(layer0_N411_wire), .M1(M1[823:822]));

wire [2:0] layer0_N412_wire = {M0[489], M0[334], M0[307]};
layer0_N412 layer0_N412_inst (.M0(layer0_N412_wire), .M1(M1[825:824]));

wire [2:0] layer0_N413_wire = {M0[398], M0[217], M0[150]};
layer0_N413 layer0_N413_inst (.M0(layer0_N413_wire), .M1(M1[827:826]));

wire [2:0] layer0_N414_wire = {M0[494], M0[366], M0[180]};
layer0_N414 layer0_N414_inst (.M0(layer0_N414_wire), .M1(M1[829:828]));

wire [2:0] layer0_N415_wire = {M0[345], M0[141], M0[58]};
layer0_N415 layer0_N415_inst (.M0(layer0_N415_wire), .M1(M1[831:830]));

wire [2:0] layer0_N416_wire = {M0[374], M0[230], M0[50]};
layer0_N416 layer0_N416_inst (.M0(layer0_N416_wire), .M1(M1[833:832]));

wire [2:0] layer0_N417_wire = {M0[302], M0[276], M0[238]};
layer0_N417 layer0_N417_inst (.M0(layer0_N417_wire), .M1(M1[835:834]));

wire [2:0] layer0_N418_wire = {M0[439], M0[364], M0[128]};
layer0_N418 layer0_N418_inst (.M0(layer0_N418_wire), .M1(M1[837:836]));

wire [2:0] layer0_N419_wire = {M0[314], M0[202], M0[177]};
layer0_N419 layer0_N419_inst (.M0(layer0_N419_wire), .M1(M1[839:838]));

wire [2:0] layer0_N420_wire = {M0[481], M0[388], M0[103]};
layer0_N420 layer0_N420_inst (.M0(layer0_N420_wire), .M1(M1[841:840]));

wire [2:0] layer0_N421_wire = {M0[470], M0[420], M0[319]};
layer0_N421 layer0_N421_inst (.M0(layer0_N421_wire), .M1(M1[843:842]));

wire [2:0] layer0_N422_wire = {M0[421], M0[294], M0[176]};
layer0_N422 layer0_N422_inst (.M0(layer0_N422_wire), .M1(M1[845:844]));

wire [2:0] layer0_N423_wire = {M0[336], M0[140], M0[90]};
layer0_N423 layer0_N423_inst (.M0(layer0_N423_wire), .M1(M1[847:846]));

wire [2:0] layer0_N424_wire = {M0[386], M0[232], M0[125]};
layer0_N424 layer0_N424_inst (.M0(layer0_N424_wire), .M1(M1[849:848]));

wire [2:0] layer0_N425_wire = {M0[490], M0[224], M0[191]};
layer0_N425 layer0_N425_inst (.M0(layer0_N425_wire), .M1(M1[851:850]));

wire [2:0] layer0_N426_wire = {M0[500], M0[287], M0[267]};
layer0_N426 layer0_N426_inst (.M0(layer0_N426_wire), .M1(M1[853:852]));

wire [2:0] layer0_N427_wire = {M0[154], M0[153], M0[132]};
layer0_N427 layer0_N427_inst (.M0(layer0_N427_wire), .M1(M1[855:854]));

wire [2:0] layer0_N428_wire = {M0[450], M0[114], M0[65]};
layer0_N428 layer0_N428_inst (.M0(layer0_N428_wire), .M1(M1[857:856]));

wire [2:0] layer0_N429_wire = {M0[340], M0[207], M0[94]};
layer0_N429 layer0_N429_inst (.M0(layer0_N429_wire), .M1(M1[859:858]));

wire [2:0] layer0_N430_wire = {M0[299], M0[288], M0[82]};
layer0_N430 layer0_N430_inst (.M0(layer0_N430_wire), .M1(M1[861:860]));

wire [2:0] layer0_N431_wire = {M0[462], M0[204], M0[107]};
layer0_N431 layer0_N431_inst (.M0(layer0_N431_wire), .M1(M1[863:862]));

wire [2:0] layer0_N432_wire = {M0[480], M0[104], M0[78]};
layer0_N432 layer0_N432_inst (.M0(layer0_N432_wire), .M1(M1[865:864]));

wire [2:0] layer0_N433_wire = {M0[240], M0[180], M0[8]};
layer0_N433 layer0_N433_inst (.M0(layer0_N433_wire), .M1(M1[867:866]));

wire [2:0] layer0_N434_wire = {M0[202], M0[199], M0[127]};
layer0_N434 layer0_N434_inst (.M0(layer0_N434_wire), .M1(M1[869:868]));

wire [2:0] layer0_N435_wire = {M0[479], M0[450], M0[124]};
layer0_N435 layer0_N435_inst (.M0(layer0_N435_wire), .M1(M1[871:870]));

wire [2:0] layer0_N436_wire = {M0[425], M0[132], M0[91]};
layer0_N436 layer0_N436_inst (.M0(layer0_N436_wire), .M1(M1[873:872]));

wire [2:0] layer0_N437_wire = {M0[470], M0[307], M0[121]};
layer0_N437 layer0_N437_inst (.M0(layer0_N437_wire), .M1(M1[875:874]));

wire [2:0] layer0_N438_wire = {M0[330], M0[195], M0[49]};
layer0_N438 layer0_N438_inst (.M0(layer0_N438_wire), .M1(M1[877:876]));

wire [2:0] layer0_N439_wire = {M0[365], M0[326], M0[161]};
layer0_N439 layer0_N439_inst (.M0(layer0_N439_wire), .M1(M1[879:878]));

wire [2:0] layer0_N440_wire = {M0[205], M0[187], M0[172]};
layer0_N440 layer0_N440_inst (.M0(layer0_N440_wire), .M1(M1[881:880]));

wire [2:0] layer0_N441_wire = {M0[257], M0[229], M0[156]};
layer0_N441 layer0_N441_inst (.M0(layer0_N441_wire), .M1(M1[883:882]));

wire [2:0] layer0_N442_wire = {M0[490], M0[378], M0[173]};
layer0_N442 layer0_N442_inst (.M0(layer0_N442_wire), .M1(M1[885:884]));

wire [2:0] layer0_N443_wire = {M0[480], M0[374], M0[280]};
layer0_N443 layer0_N443_inst (.M0(layer0_N443_wire), .M1(M1[887:886]));

wire [2:0] layer0_N444_wire = {M0[285], M0[270], M0[30]};
layer0_N444 layer0_N444_inst (.M0(layer0_N444_wire), .M1(M1[889:888]));

wire [2:0] layer0_N445_wire = {M0[406], M0[389], M0[357]};
layer0_N445 layer0_N445_inst (.M0(layer0_N445_wire), .M1(M1[891:890]));

wire [2:0] layer0_N446_wire = {M0[390], M0[92], M0[67]};
layer0_N446 layer0_N446_inst (.M0(layer0_N446_wire), .M1(M1[893:892]));

wire [2:0] layer0_N447_wire = {M0[420], M0[311], M0[102]};
layer0_N447 layer0_N447_inst (.M0(layer0_N447_wire), .M1(M1[895:894]));

wire [2:0] layer0_N448_wire = {M0[312], M0[220], M0[214]};
layer0_N448 layer0_N448_inst (.M0(layer0_N448_wire), .M1(M1[897:896]));

wire [2:0] layer0_N449_wire = {M0[290], M0[172], M0[17]};
layer0_N449 layer0_N449_inst (.M0(layer0_N449_wire), .M1(M1[899:898]));

wire [2:0] layer0_N450_wire = {M0[366], M0[295], M0[242]};
layer0_N450 layer0_N450_inst (.M0(layer0_N450_wire), .M1(M1[901:900]));

wire [2:0] layer0_N451_wire = {M0[466], M0[346], M0[230]};
layer0_N451 layer0_N451_inst (.M0(layer0_N451_wire), .M1(M1[903:902]));

wire [2:0] layer0_N452_wire = {M0[380], M0[321], M0[149]};
layer0_N452 layer0_N452_inst (.M0(layer0_N452_wire), .M1(M1[905:904]));

wire [2:0] layer0_N453_wire = {M0[215], M0[144], M0[8]};
layer0_N453 layer0_N453_inst (.M0(layer0_N453_wire), .M1(M1[907:906]));

wire [2:0] layer0_N454_wire = {M0[191], M0[188], M0[5]};
layer0_N454 layer0_N454_inst (.M0(layer0_N454_wire), .M1(M1[909:908]));

wire [2:0] layer0_N455_wire = {M0[104], M0[80], M0[23]};
layer0_N455 layer0_N455_inst (.M0(layer0_N455_wire), .M1(M1[911:910]));

wire [2:0] layer0_N456_wire = {M0[334], M0[314], M0[72]};
layer0_N456 layer0_N456_inst (.M0(layer0_N456_wire), .M1(M1[913:912]));

wire [2:0] layer0_N457_wire = {M0[431], M0[249], M0[198]};
layer0_N457 layer0_N457_inst (.M0(layer0_N457_wire), .M1(M1[915:914]));

wire [2:0] layer0_N458_wire = {M0[390], M0[357], M0[173]};
layer0_N458 layer0_N458_inst (.M0(layer0_N458_wire), .M1(M1[917:916]));

wire [2:0] layer0_N459_wire = {M0[137], M0[97], M0[91]};
layer0_N459 layer0_N459_inst (.M0(layer0_N459_wire), .M1(M1[919:918]));

wire [2:0] layer0_N460_wire = {M0[471], M0[100], M0[17]};
layer0_N460 layer0_N460_inst (.M0(layer0_N460_wire), .M1(M1[921:920]));

wire [2:0] layer0_N461_wire = {M0[399], M0[250], M0[10]};
layer0_N461 layer0_N461_inst (.M0(layer0_N461_wire), .M1(M1[923:922]));

wire [2:0] layer0_N462_wire = {M0[428], M0[356], M0[243]};
layer0_N462 layer0_N462_inst (.M0(layer0_N462_wire), .M1(M1[925:924]));

wire [2:0] layer0_N463_wire = {M0[454], M0[315], M0[102]};
layer0_N463 layer0_N463_inst (.M0(layer0_N463_wire), .M1(M1[927:926]));

wire [2:0] layer0_N464_wire = {M0[484], M0[256], M0[190]};
layer0_N464 layer0_N464_inst (.M0(layer0_N464_wire), .M1(M1[929:928]));

wire [2:0] layer0_N465_wire = {M0[366], M0[127], M0[19]};
layer0_N465 layer0_N465_inst (.M0(layer0_N465_wire), .M1(M1[931:930]));

wire [2:0] layer0_N466_wire = {M0[293], M0[247], M0[125]};
layer0_N466 layer0_N466_inst (.M0(layer0_N466_wire), .M1(M1[933:932]));

wire [2:0] layer0_N467_wire = {M0[296], M0[88], M0[47]};
layer0_N467 layer0_N467_inst (.M0(layer0_N467_wire), .M1(M1[935:934]));

wire [2:0] layer0_N468_wire = {M0[480], M0[448], M0[216]};
layer0_N468 layer0_N468_inst (.M0(layer0_N468_wire), .M1(M1[937:936]));

wire [2:0] layer0_N469_wire = {M0[433], M0[153], M0[25]};
layer0_N469 layer0_N469_inst (.M0(layer0_N469_wire), .M1(M1[939:938]));

wire [2:0] layer0_N470_wire = {M0[419], M0[125], M0[57]};
layer0_N470 layer0_N470_inst (.M0(layer0_N470_wire), .M1(M1[941:940]));

wire [2:0] layer0_N471_wire = {M0[262], M0[96], M0[71]};
layer0_N471 layer0_N471_inst (.M0(layer0_N471_wire), .M1(M1[943:942]));

wire [2:0] layer0_N472_wire = {M0[352], M0[208], M0[64]};
layer0_N472 layer0_N472_inst (.M0(layer0_N472_wire), .M1(M1[945:944]));

wire [2:0] layer0_N473_wire = {M0[134], M0[98], M0[16]};
layer0_N473 layer0_N473_inst (.M0(layer0_N473_wire), .M1(M1[947:946]));

wire [2:0] layer0_N474_wire = {M0[506], M0[333], M0[206]};
layer0_N474 layer0_N474_inst (.M0(layer0_N474_wire), .M1(M1[949:948]));

wire [2:0] layer0_N475_wire = {M0[431], M0[416], M0[383]};
layer0_N475 layer0_N475_inst (.M0(layer0_N475_wire), .M1(M1[951:950]));

wire [2:0] layer0_N476_wire = {M0[466], M0[128], M0[25]};
layer0_N476 layer0_N476_inst (.M0(layer0_N476_wire), .M1(M1[953:952]));

wire [2:0] layer0_N477_wire = {M0[336], M0[164], M0[75]};
layer0_N477 layer0_N477_inst (.M0(layer0_N477_wire), .M1(M1[955:954]));

wire [2:0] layer0_N478_wire = {M0[285], M0[141], M0[12]};
layer0_N478 layer0_N478_inst (.M0(layer0_N478_wire), .M1(M1[957:956]));

wire [2:0] layer0_N479_wire = {M0[253], M0[100], M0[7]};
layer0_N479 layer0_N479_inst (.M0(layer0_N479_wire), .M1(M1[959:958]));

wire [2:0] layer0_N480_wire = {M0[299], M0[121], M0[46]};
layer0_N480 layer0_N480_inst (.M0(layer0_N480_wire), .M1(M1[961:960]));

wire [2:0] layer0_N481_wire = {M0[279], M0[224], M0[47]};
layer0_N481 layer0_N481_inst (.M0(layer0_N481_wire), .M1(M1[963:962]));

wire [2:0] layer0_N482_wire = {M0[363], M0[192], M0[45]};
layer0_N482 layer0_N482_inst (.M0(layer0_N482_wire), .M1(M1[965:964]));

wire [2:0] layer0_N483_wire = {M0[478], M0[316], M0[98]};
layer0_N483 layer0_N483_inst (.M0(layer0_N483_wire), .M1(M1[967:966]));

wire [2:0] layer0_N484_wire = {M0[374], M0[214], M0[73]};
layer0_N484 layer0_N484_inst (.M0(layer0_N484_wire), .M1(M1[969:968]));

wire [2:0] layer0_N485_wire = {M0[448], M0[349], M0[334]};
layer0_N485 layer0_N485_inst (.M0(layer0_N485_wire), .M1(M1[971:970]));

wire [2:0] layer0_N486_wire = {M0[476], M0[171], M0[134]};
layer0_N486 layer0_N486_inst (.M0(layer0_N486_wire), .M1(M1[973:972]));

wire [2:0] layer0_N487_wire = {M0[363], M0[282], M0[86]};
layer0_N487 layer0_N487_inst (.M0(layer0_N487_wire), .M1(M1[975:974]));

wire [2:0] layer0_N488_wire = {M0[348], M0[260], M0[6]};
layer0_N488 layer0_N488_inst (.M0(layer0_N488_wire), .M1(M1[977:976]));

wire [2:0] layer0_N489_wire = {M0[443], M0[153], M0[131]};
layer0_N489 layer0_N489_inst (.M0(layer0_N489_wire), .M1(M1[979:978]));

wire [2:0] layer0_N490_wire = {M0[132], M0[95], M0[50]};
layer0_N490 layer0_N490_inst (.M0(layer0_N490_wire), .M1(M1[981:980]));

wire [2:0] layer0_N491_wire = {M0[455], M0[408], M0[176]};
layer0_N491 layer0_N491_inst (.M0(layer0_N491_wire), .M1(M1[983:982]));

wire [2:0] layer0_N492_wire = {M0[476], M0[307], M0[18]};
layer0_N492 layer0_N492_inst (.M0(layer0_N492_wire), .M1(M1[985:984]));

wire [2:0] layer0_N493_wire = {M0[449], M0[269], M0[145]};
layer0_N493 layer0_N493_inst (.M0(layer0_N493_wire), .M1(M1[987:986]));

wire [2:0] layer0_N494_wire = {M0[491], M0[370], M0[103]};
layer0_N494 layer0_N494_inst (.M0(layer0_N494_wire), .M1(M1[989:988]));

wire [2:0] layer0_N495_wire = {M0[468], M0[330], M0[141]};
layer0_N495 layer0_N495_inst (.M0(layer0_N495_wire), .M1(M1[991:990]));

wire [2:0] layer0_N496_wire = {M0[406], M0[115], M0[5]};
layer0_N496 layer0_N496_inst (.M0(layer0_N496_wire), .M1(M1[993:992]));

wire [2:0] layer0_N497_wire = {M0[388], M0[329], M0[242]};
layer0_N497 layer0_N497_inst (.M0(layer0_N497_wire), .M1(M1[995:994]));

wire [2:0] layer0_N498_wire = {M0[401], M0[172], M0[122]};
layer0_N498 layer0_N498_inst (.M0(layer0_N498_wire), .M1(M1[997:996]));

wire [2:0] layer0_N499_wire = {M0[461], M0[265], M0[152]};
layer0_N499 layer0_N499_inst (.M0(layer0_N499_wire), .M1(M1[999:998]));

wire [2:0] layer0_N500_wire = {M0[502], M0[354], M0[186]};
layer0_N500 layer0_N500_inst (.M0(layer0_N500_wire), .M1(M1[1001:1000]));

wire [2:0] layer0_N501_wire = {M0[442], M0[398], M0[103]};
layer0_N501 layer0_N501_inst (.M0(layer0_N501_wire), .M1(M1[1003:1002]));

wire [2:0] layer0_N502_wire = {M0[442], M0[249], M0[68]};
layer0_N502 layer0_N502_inst (.M0(layer0_N502_wire), .M1(M1[1005:1004]));

wire [2:0] layer0_N503_wire = {M0[249], M0[199], M0[87]};
layer0_N503 layer0_N503_inst (.M0(layer0_N503_wire), .M1(M1[1007:1006]));

wire [2:0] layer0_N504_wire = {M0[400], M0[390], M0[389]};
layer0_N504 layer0_N504_inst (.M0(layer0_N504_wire), .M1(M1[1009:1008]));

wire [2:0] layer0_N505_wire = {M0[249], M0[191], M0[71]};
layer0_N505 layer0_N505_inst (.M0(layer0_N505_wire), .M1(M1[1011:1010]));

wire [2:0] layer0_N506_wire = {M0[505], M0[284], M0[185]};
layer0_N506 layer0_N506_inst (.M0(layer0_N506_wire), .M1(M1[1013:1012]));

wire [2:0] layer0_N507_wire = {M0[490], M0[179], M0[11]};
layer0_N507 layer0_N507_inst (.M0(layer0_N507_wire), .M1(M1[1015:1014]));

wire [2:0] layer0_N508_wire = {M0[429], M0[99], M0[36]};
layer0_N508 layer0_N508_inst (.M0(layer0_N508_wire), .M1(M1[1017:1016]));

wire [2:0] layer0_N509_wire = {M0[369], M0[95], M0[14]};
layer0_N509 layer0_N509_inst (.M0(layer0_N509_wire), .M1(M1[1019:1018]));

wire [2:0] layer0_N510_wire = {M0[467], M0[443], M0[139]};
layer0_N510 layer0_N510_inst (.M0(layer0_N510_wire), .M1(M1[1021:1020]));

wire [2:0] layer0_N511_wire = {M0[262], M0[76], M0[54]};
layer0_N511 layer0_N511_inst (.M0(layer0_N511_wire), .M1(M1[1023:1022]));

wire [2:0] layer0_N512_wire = {M0[510], M0[396], M0[308]};
layer0_N512 layer0_N512_inst (.M0(layer0_N512_wire), .M1(M1[1025:1024]));

wire [2:0] layer0_N513_wire = {M0[211], M0[150], M0[13]};
layer0_N513 layer0_N513_inst (.M0(layer0_N513_wire), .M1(M1[1027:1026]));

wire [2:0] layer0_N514_wire = {M0[456], M0[101], M0[75]};
layer0_N514 layer0_N514_inst (.M0(layer0_N514_wire), .M1(M1[1029:1028]));

wire [2:0] layer0_N515_wire = {M0[287], M0[179], M0[103]};
layer0_N515 layer0_N515_inst (.M0(layer0_N515_wire), .M1(M1[1031:1030]));

wire [2:0] layer0_N516_wire = {M0[443], M0[343], M0[268]};
layer0_N516 layer0_N516_inst (.M0(layer0_N516_wire), .M1(M1[1033:1032]));

wire [2:0] layer0_N517_wire = {M0[493], M0[120], M0[50]};
layer0_N517 layer0_N517_inst (.M0(layer0_N517_wire), .M1(M1[1035:1034]));

wire [2:0] layer0_N518_wire = {M0[510], M0[405], M0[37]};
layer0_N518 layer0_N518_inst (.M0(layer0_N518_wire), .M1(M1[1037:1036]));

wire [2:0] layer0_N519_wire = {M0[90], M0[51], M0[4]};
layer0_N519 layer0_N519_inst (.M0(layer0_N519_wire), .M1(M1[1039:1038]));

wire [2:0] layer0_N520_wire = {M0[319], M0[257], M0[232]};
layer0_N520 layer0_N520_inst (.M0(layer0_N520_wire), .M1(M1[1041:1040]));

wire [2:0] layer0_N521_wire = {M0[504], M0[452], M0[202]};
layer0_N521 layer0_N521_inst (.M0(layer0_N521_wire), .M1(M1[1043:1042]));

wire [2:0] layer0_N522_wire = {M0[428], M0[354], M0[136]};
layer0_N522 layer0_N522_inst (.M0(layer0_N522_wire), .M1(M1[1045:1044]));

wire [2:0] layer0_N523_wire = {M0[370], M0[244], M0[85]};
layer0_N523 layer0_N523_inst (.M0(layer0_N523_wire), .M1(M1[1047:1046]));

wire [2:0] layer0_N524_wire = {M0[276], M0[105], M0[97]};
layer0_N524 layer0_N524_inst (.M0(layer0_N524_wire), .M1(M1[1049:1048]));

wire [2:0] layer0_N525_wire = {M0[442], M0[265], M0[251]};
layer0_N525 layer0_N525_inst (.M0(layer0_N525_wire), .M1(M1[1051:1050]));

wire [2:0] layer0_N526_wire = {M0[434], M0[82], M0[3]};
layer0_N526 layer0_N526_inst (.M0(layer0_N526_wire), .M1(M1[1053:1052]));

wire [2:0] layer0_N527_wire = {M0[397], M0[281], M0[117]};
layer0_N527 layer0_N527_inst (.M0(layer0_N527_wire), .M1(M1[1055:1054]));

wire [2:0] layer0_N528_wire = {M0[447], M0[76], M0[1]};
layer0_N528 layer0_N528_inst (.M0(layer0_N528_wire), .M1(M1[1057:1056]));

wire [2:0] layer0_N529_wire = {M0[505], M0[455], M0[397]};
layer0_N529 layer0_N529_inst (.M0(layer0_N529_wire), .M1(M1[1059:1058]));

wire [2:0] layer0_N530_wire = {M0[341], M0[324], M0[146]};
layer0_N530 layer0_N530_inst (.M0(layer0_N530_wire), .M1(M1[1061:1060]));

wire [2:0] layer0_N531_wire = {M0[490], M0[332], M0[78]};
layer0_N531 layer0_N531_inst (.M0(layer0_N531_wire), .M1(M1[1063:1062]));

wire [2:0] layer0_N532_wire = {M0[477], M0[102], M0[76]};
layer0_N532 layer0_N532_inst (.M0(layer0_N532_wire), .M1(M1[1065:1064]));

wire [2:0] layer0_N533_wire = {M0[489], M0[195], M0[73]};
layer0_N533 layer0_N533_inst (.M0(layer0_N533_wire), .M1(M1[1067:1066]));

wire [2:0] layer0_N534_wire = {M0[271], M0[177], M0[44]};
layer0_N534 layer0_N534_inst (.M0(layer0_N534_wire), .M1(M1[1069:1068]));

wire [2:0] layer0_N535_wire = {M0[427], M0[365], M0[265]};
layer0_N535 layer0_N535_inst (.M0(layer0_N535_wire), .M1(M1[1071:1070]));

wire [2:0] layer0_N536_wire = {M0[125], M0[46], M0[24]};
layer0_N536 layer0_N536_inst (.M0(layer0_N536_wire), .M1(M1[1073:1072]));

wire [2:0] layer0_N537_wire = {M0[351], M0[101], M0[84]};
layer0_N537 layer0_N537_inst (.M0(layer0_N537_wire), .M1(M1[1075:1074]));

wire [2:0] layer0_N538_wire = {M0[374], M0[312], M0[94]};
layer0_N538 layer0_N538_inst (.M0(layer0_N538_wire), .M1(M1[1077:1076]));

wire [2:0] layer0_N539_wire = {M0[352], M0[332], M0[146]};
layer0_N539 layer0_N539_inst (.M0(layer0_N539_wire), .M1(M1[1079:1078]));

wire [2:0] layer0_N540_wire = {M0[504], M0[454], M0[179]};
layer0_N540 layer0_N540_inst (.M0(layer0_N540_wire), .M1(M1[1081:1080]));

wire [2:0] layer0_N541_wire = {M0[373], M0[370], M0[248]};
layer0_N541 layer0_N541_inst (.M0(layer0_N541_wire), .M1(M1[1083:1082]));

wire [2:0] layer0_N542_wire = {M0[259], M0[231], M0[105]};
layer0_N542 layer0_N542_inst (.M0(layer0_N542_wire), .M1(M1[1085:1084]));

wire [2:0] layer0_N543_wire = {M0[491], M0[467], M0[19]};
layer0_N543 layer0_N543_inst (.M0(layer0_N543_wire), .M1(M1[1087:1086]));

wire [2:0] layer0_N544_wire = {M0[490], M0[196], M0[137]};
layer0_N544 layer0_N544_inst (.M0(layer0_N544_wire), .M1(M1[1089:1088]));

wire [2:0] layer0_N545_wire = {M0[382], M0[292], M0[252]};
layer0_N545 layer0_N545_inst (.M0(layer0_N545_wire), .M1(M1[1091:1090]));

wire [2:0] layer0_N546_wire = {M0[447], M0[350], M0[78]};
layer0_N546 layer0_N546_inst (.M0(layer0_N546_wire), .M1(M1[1093:1092]));

wire [2:0] layer0_N547_wire = {M0[285], M0[119], M0[38]};
layer0_N547 layer0_N547_inst (.M0(layer0_N547_wire), .M1(M1[1095:1094]));

wire [2:0] layer0_N548_wire = {M0[457], M0[389], M0[184]};
layer0_N548 layer0_N548_inst (.M0(layer0_N548_wire), .M1(M1[1097:1096]));

wire [2:0] layer0_N549_wire = {M0[485], M0[365], M0[224]};
layer0_N549 layer0_N549_inst (.M0(layer0_N549_wire), .M1(M1[1099:1098]));

wire [2:0] layer0_N550_wire = {M0[498], M0[29], M0[8]};
layer0_N550 layer0_N550_inst (.M0(layer0_N550_wire), .M1(M1[1101:1100]));

wire [2:0] layer0_N551_wire = {M0[510], M0[219], M0[113]};
layer0_N551 layer0_N551_inst (.M0(layer0_N551_wire), .M1(M1[1103:1102]));

wire [2:0] layer0_N552_wire = {M0[317], M0[285], M0[58]};
layer0_N552 layer0_N552_inst (.M0(layer0_N552_wire), .M1(M1[1105:1104]));

wire [2:0] layer0_N553_wire = {M0[482], M0[256], M0[38]};
layer0_N553 layer0_N553_inst (.M0(layer0_N553_wire), .M1(M1[1107:1106]));

wire [2:0] layer0_N554_wire = {M0[307], M0[306], M0[261]};
layer0_N554 layer0_N554_inst (.M0(layer0_N554_wire), .M1(M1[1109:1108]));

wire [2:0] layer0_N555_wire = {M0[468], M0[351], M0[162]};
layer0_N555 layer0_N555_inst (.M0(layer0_N555_wire), .M1(M1[1111:1110]));

wire [2:0] layer0_N556_wire = {M0[459], M0[403], M0[243]};
layer0_N556 layer0_N556_inst (.M0(layer0_N556_wire), .M1(M1[1113:1112]));

wire [2:0] layer0_N557_wire = {M0[481], M0[389], M0[275]};
layer0_N557 layer0_N557_inst (.M0(layer0_N557_wire), .M1(M1[1115:1114]));

wire [2:0] layer0_N558_wire = {M0[488], M0[169], M0[81]};
layer0_N558 layer0_N558_inst (.M0(layer0_N558_wire), .M1(M1[1117:1116]));

wire [2:0] layer0_N559_wire = {M0[309], M0[246], M0[16]};
layer0_N559 layer0_N559_inst (.M0(layer0_N559_wire), .M1(M1[1119:1118]));

wire [2:0] layer0_N560_wire = {M0[396], M0[337], M0[50]};
layer0_N560 layer0_N560_inst (.M0(layer0_N560_wire), .M1(M1[1121:1120]));

wire [2:0] layer0_N561_wire = {M0[486], M0[219], M0[112]};
layer0_N561 layer0_N561_inst (.M0(layer0_N561_wire), .M1(M1[1123:1122]));

wire [2:0] layer0_N562_wire = {M0[424], M0[181], M0[160]};
layer0_N562 layer0_N562_inst (.M0(layer0_N562_wire), .M1(M1[1125:1124]));

wire [2:0] layer0_N563_wire = {M0[401], M0[94], M0[65]};
layer0_N563 layer0_N563_inst (.M0(layer0_N563_wire), .M1(M1[1127:1126]));

wire [2:0] layer0_N564_wire = {M0[509], M0[282], M0[228]};
layer0_N564 layer0_N564_inst (.M0(layer0_N564_wire), .M1(M1[1129:1128]));

wire [2:0] layer0_N565_wire = {M0[369], M0[261], M0[105]};
layer0_N565 layer0_N565_inst (.M0(layer0_N565_wire), .M1(M1[1131:1130]));

wire [2:0] layer0_N566_wire = {M0[285], M0[206], M0[95]};
layer0_N566 layer0_N566_inst (.M0(layer0_N566_wire), .M1(M1[1133:1132]));

wire [2:0] layer0_N567_wire = {M0[392], M0[360], M0[264]};
layer0_N567 layer0_N567_inst (.M0(layer0_N567_wire), .M1(M1[1135:1134]));

wire [2:0] layer0_N568_wire = {M0[486], M0[81], M0[75]};
layer0_N568 layer0_N568_inst (.M0(layer0_N568_wire), .M1(M1[1137:1136]));

wire [2:0] layer0_N569_wire = {M0[480], M0[209], M0[118]};
layer0_N569 layer0_N569_inst (.M0(layer0_N569_wire), .M1(M1[1139:1138]));

wire [2:0] layer0_N570_wire = {M0[237], M0[174], M0[115]};
layer0_N570 layer0_N570_inst (.M0(layer0_N570_wire), .M1(M1[1141:1140]));

wire [2:0] layer0_N571_wire = {M0[232], M0[101], M0[84]};
layer0_N571 layer0_N571_inst (.M0(layer0_N571_wire), .M1(M1[1143:1142]));

wire [2:0] layer0_N572_wire = {M0[500], M0[331], M0[240]};
layer0_N572 layer0_N572_inst (.M0(layer0_N572_wire), .M1(M1[1145:1144]));

wire [2:0] layer0_N573_wire = {M0[329], M0[167], M0[16]};
layer0_N573 layer0_N573_inst (.M0(layer0_N573_wire), .M1(M1[1147:1146]));

wire [2:0] layer0_N574_wire = {M0[420], M0[252], M0[108]};
layer0_N574 layer0_N574_inst (.M0(layer0_N574_wire), .M1(M1[1149:1148]));

wire [2:0] layer0_N575_wire = {M0[176], M0[79], M0[69]};
layer0_N575 layer0_N575_inst (.M0(layer0_N575_wire), .M1(M1[1151:1150]));

wire [2:0] layer0_N576_wire = {M0[478], M0[472], M0[374]};
layer0_N576 layer0_N576_inst (.M0(layer0_N576_wire), .M1(M1[1153:1152]));

wire [2:0] layer0_N577_wire = {M0[508], M0[219], M0[165]};
layer0_N577 layer0_N577_inst (.M0(layer0_N577_wire), .M1(M1[1155:1154]));

wire [2:0] layer0_N578_wire = {M0[483], M0[342], M0[251]};
layer0_N578 layer0_N578_inst (.M0(layer0_N578_wire), .M1(M1[1157:1156]));

wire [2:0] layer0_N579_wire = {M0[328], M0[196], M0[150]};
layer0_N579 layer0_N579_inst (.M0(layer0_N579_wire), .M1(M1[1159:1158]));

wire [2:0] layer0_N580_wire = {M0[477], M0[422], M0[76]};
layer0_N580 layer0_N580_inst (.M0(layer0_N580_wire), .M1(M1[1161:1160]));

wire [2:0] layer0_N581_wire = {M0[177], M0[73], M0[66]};
layer0_N581 layer0_N581_inst (.M0(layer0_N581_wire), .M1(M1[1163:1162]));

wire [2:0] layer0_N582_wire = {M0[344], M0[264], M0[35]};
layer0_N582 layer0_N582_inst (.M0(layer0_N582_wire), .M1(M1[1165:1164]));

wire [2:0] layer0_N583_wire = {M0[340], M0[104], M0[88]};
layer0_N583 layer0_N583_inst (.M0(layer0_N583_wire), .M1(M1[1167:1166]));

wire [2:0] layer0_N584_wire = {M0[250], M0[62], M0[40]};
layer0_N584 layer0_N584_inst (.M0(layer0_N584_wire), .M1(M1[1169:1168]));

wire [2:0] layer0_N585_wire = {M0[434], M0[421], M0[51]};
layer0_N585 layer0_N585_inst (.M0(layer0_N585_wire), .M1(M1[1171:1170]));

wire [2:0] layer0_N586_wire = {M0[73], M0[41], M0[38]};
layer0_N586 layer0_N586_inst (.M0(layer0_N586_wire), .M1(M1[1173:1172]));

wire [2:0] layer0_N587_wire = {M0[391], M0[321], M0[39]};
layer0_N587 layer0_N587_inst (.M0(layer0_N587_wire), .M1(M1[1175:1174]));

wire [2:0] layer0_N588_wire = {M0[109], M0[63], M0[24]};
layer0_N588 layer0_N588_inst (.M0(layer0_N588_wire), .M1(M1[1177:1176]));

wire [2:0] layer0_N589_wire = {M0[451], M0[233], M0[212]};
layer0_N589 layer0_N589_inst (.M0(layer0_N589_wire), .M1(M1[1179:1178]));

wire [2:0] layer0_N590_wire = {M0[501], M0[241], M0[110]};
layer0_N590 layer0_N590_inst (.M0(layer0_N590_wire), .M1(M1[1181:1180]));

wire [2:0] layer0_N591_wire = {M0[401], M0[339], M0[238]};
layer0_N591 layer0_N591_inst (.M0(layer0_N591_wire), .M1(M1[1183:1182]));

wire [2:0] layer0_N592_wire = {M0[330], M0[148], M0[63]};
layer0_N592 layer0_N592_inst (.M0(layer0_N592_wire), .M1(M1[1185:1184]));

endmodule